module rams_sp_rom0_8_sec (clk, enA, enB, addrA, addrB, doA, doB);
input clk;
input enA, enB;
input [11:0] addrA, addrB;
output [31:0] doA, doB;
(*rom_style = "block" *) reg [2751:0] dataA, dataB;
always @(posedge clk)
begin
if (enA)
case(addrA)
12'b000000000000: dataA <= 32'b11100101001110101110000110111000;
12'b000000000001: dataA <= 32'b00001000100111101110010000011101;
12'b000000000010: dataA <= 32'b01001000011001011011100010101110;
12'b000000000011: dataA <= 32'b00000011100011010110001100110001;
12'b000000000100: dataA <= 32'b01010100110010110111011011110110;
12'b000000000101: dataA <= 32'b00000101100001100000001001111011;
12'b000000000110: dataA <= 32'b01001011101000111011000001001011;
12'b000000000111: dataA <= 32'b00001000110100101111001101010111;
12'b000000001000: dataA <= 32'b11110100010100101011111101001100;
12'b000000001001: dataA <= 32'b00000110001011100100100011001001;
12'b000000001010: dataA <= 32'b00100001000001111101110101010101;
12'b000000001011: dataA <= 32'b00000010111010110111011101011101;
12'b000000001100: dataA <= 32'b10110111001000101010100101001000;
12'b000000001101: dataA <= 32'b00000001110010010001000011101101;
12'b000000001110: dataA <= 32'b00110000111110111110011110110101;
12'b000000001111: dataA <= 32'b00000011111011010111011110011100;
12'b000000010000: dataA <= 32'b10101100001001101111100100011010;
12'b000000010001: dataA <= 32'b00000101101000011100001100010010;
12'b000000010010: dataA <= 32'b11011001001010110101000011010011;
12'b000000010011: dataA <= 32'b00001001100010011100001100110100;
12'b000000010100: dataA <= 32'b01011100011111000111000011010110;
12'b000000010101: dataA <= 32'b00001111001110010100111001001010;
12'b000000010110: dataA <= 32'b10110011000101000011110110101101;
12'b000000010111: dataA <= 32'b00000001001100000110011100101101;
12'b000000011000: dataA <= 32'b00001100010010101001100100100111;
12'b000000011001: dataA <= 32'b00000111011110100101100101011010;
12'b000000011010: dataA <= 32'b10101010100010011111100111110111;
12'b000000011011: dataA <= 32'b00001001100001110000001110000010;
12'b000000011100: dataA <= 32'b10010101001011011110010110110001;
12'b000000011101: dataA <= 32'b00000001001111100100101110000100;
12'b000000011110: dataA <= 32'b10001100111110110111011000111000;
12'b000000011111: dataA <= 32'b00001001100101001000011010010011;
12'b000000100000: dataA <= 32'b01000011001111010101000001110110;
12'b000000100001: dataA <= 32'b00000101010100110001001010011100;
12'b000000100010: dataA <= 32'b10111100111101001011001101100101;
12'b000000100011: dataA <= 32'b00000110010111001111011001000100;
12'b000000100100: dataA <= 32'b10010010010110011110001100010110;
12'b000000100101: dataA <= 32'b00001100101010110010010001011010;
12'b000000100110: dataA <= 32'b11110110011000101101110101010100;
12'b000000100111: dataA <= 32'b00001011110101011101010010110001;
12'b000000101000: dataA <= 32'b11000100110000111010000001001000;
12'b000000101001: dataA <= 32'b00000010011001010001100001101010;
12'b000000101010: dataA <= 32'b00010111101101011011111000001101;
12'b000000101011: dataA <= 32'b00001001101001001110001101000111;
12'b000000101100: dataA <= 32'b00101100111100010011001110000111;
12'b000000101101: dataA <= 32'b00001011110000100010111011110100;
12'b000000101110: dataA <= 32'b10010000110001100011011100001010;
12'b000000101111: dataA <= 32'b00001000010111101011010100001011;
12'b000000110000: dataA <= 32'b11011010111001100110001000110011;
12'b000000110001: dataA <= 32'b00001101111001000011001100011100;
12'b000000110010: dataA <= 32'b00101011011010000011100001001110;
12'b000000110011: dataA <= 32'b00000100110101011101010001000111;
12'b000000110100: dataA <= 32'b01110100011010000010000101101001;
12'b000000110101: dataA <= 32'b00000011100011101000001000111010;
12'b000000110110: dataA <= 32'b01000011001101000110010110111000;
12'b000000110111: dataA <= 32'b00001001000101011000010111000100;
12'b000000111000: dataA <= 32'b11001110111111110011010001001111;
12'b000000111001: dataA <= 32'b00000100100010001010010111000011;
12'b000000111010: dataA <= 32'b01101010101101111011000001001000;
12'b000000111011: dataA <= 32'b00000100001110111100101000101011;
12'b000000111100: dataA <= 32'b10010111011110110111011101111001;
12'b000000111101: dataA <= 32'b00001011001111111100110101111111;
12'b000000111110: dataA <= 32'b10101000011100111010100110101001;
12'b000000111111: dataA <= 32'b00001010001011011100101100110010;
12'b000001000000: dataA <= 32'b10010001010101111110101110110110;
12'b000001000001: dataA <= 32'b00000001110010110100110101000110;
12'b000001000010: dataA <= 32'b11000111001101011110100010111001;
12'b000001000011: dataA <= 32'b00000100111101000111100001010100;
12'b000001000100: dataA <= 32'b01100010101100100110011111010001;
12'b000001000101: dataA <= 32'b00000010011001000111011001100011;
12'b000001000110: dataA <= 32'b00100101001010000010010111100001;
12'b000001000111: dataA <= 32'b00001011100101001010011101000101;
12'b000001001000: dataA <= 32'b00110001010101001110111011011001;
12'b000001001001: dataA <= 32'b00001010001001110010100000011110;
12'b000001001010: dataA <= 32'b01100101001110010001110110101000;
12'b000001001011: dataA <= 32'b00001101110001010111001011011110;
12'b000001001100: dataA <= 32'b10001011010110101011000111101101;
12'b000001001101: dataA <= 32'b00001000110001011001001011110100;
12'b000001001110: dataA <= 32'b00011111000000101110101000010101;
12'b000001001111: dataA <= 32'b00000110100111100010001010100100;
12'b000001010000: dataA <= 32'b11010010111100111100111011110001;
12'b000001010001: dataA <= 32'b00000111111011101011100001110011;
12'b000001010010: dataA <= 32'b01011100001110101100110101010011;
12'b000001010011: dataA <= 32'b00001101011011110001010010011001;
12'b000001010100: dataA <= 32'b10010011100110101111101001110110;
12'b000001010101: dataA <= 32'b00000111111110100001011001110110;
12'b000001010110: dataA <= 32'b10100111001110111101110111111000;
12'b000001010111: dataA <= 32'b00000111100111101010001000100110;
12'b000001011000: dataA <= 32'b11000100100001011011110010110000;
12'b000001011001: dataA <= 32'b00000010000101010010010000101001;
12'b000001011010: dataA <= 32'b01010100110111001110111100010100;
12'b000001011011: dataA <= 32'b00000100000010011100001001111011;
12'b000001011100: dataA <= 32'b10001111110000111011100000101110;
12'b000001011101: dataA <= 32'b00001001010100101111000101101111;
12'b000001011110: dataA <= 32'b01101110001100110100011100101010;
12'b000001011111: dataA <= 32'b00000101101100100000100010111001;
12'b000001100000: dataA <= 32'b01100001000010001101100101110110;
12'b000001100001: dataA <= 32'b00000011111100111011010101100101;
12'b000001100010: dataA <= 32'b11110111000000100011000100001001;
12'b000001100011: dataA <= 32'b00000001110100010001001011110100;
12'b000001100100: dataA <= 32'b00110000110111001101111111010010;
12'b000001100101: dataA <= 32'b00000100111101011011100010011100;
12'b000001100110: dataA <= 32'b01100110000110000111100101011100;
12'b000001100111: dataA <= 32'b00000100101001011000001100001011;
12'b000001101000: dataA <= 32'b01011001001110111100110011110101;
12'b000001101001: dataA <= 32'b00001000100010011000001100111101;
12'b000001101010: dataA <= 32'b11011000011111010110100100011000;
12'b000001101011: dataA <= 32'b00001111001011010100111101000010;
12'b000001101100: dataA <= 32'b11110010111101001100010110101101;
12'b000001101101: dataA <= 32'b00000001001110000100101000110101;
12'b000001101110: dataA <= 32'b01001000011010011001010011101001;
12'b000001101111: dataA <= 32'b00001000111110101001100001001010;
12'b000001110000: dataA <= 32'b10100110011110110111011000110110;
12'b000001110001: dataA <= 32'b00001000000001101010001001111010;
12'b000001110010: dataA <= 32'b10010101001111101101110110110001;
12'b000001110011: dataA <= 32'b00000001010001100010101110000100;
12'b000001110100: dataA <= 32'b10001111000111001110111001111000;
12'b000001110101: dataA <= 32'b00001000100100000100100010010011;
12'b000001110110: dataA <= 32'b01000101011011011100100010111000;
12'b000001110111: dataA <= 32'b00000101110101110001000010011100;
12'b000001111000: dataA <= 32'b00111100110001001011011100100100;
12'b000001111001: dataA <= 32'b00000111010111010011100001000101;
12'b000001111010: dataA <= 32'b11010000011010101101111100110100;
12'b000001111011: dataA <= 32'b00001100001000101110001101010010;
12'b000001111100: dataA <= 32'b10110010010000111110000101110101;
12'b000001111101: dataA <= 32'b00001100010011011111010010100001;
12'b000001111110: dataA <= 32'b11000100111000110010100000101011;
12'b000001111111: dataA <= 32'b00000011011011010101100101100010;
12'b000010000000: dataA <= 32'b10011011110001011100001000001101;
12'b000010000001: dataA <= 32'b00001001001001001000010101011111;
12'b000010000010: dataA <= 32'b01101100110100010011101101000100;
12'b000010000011: dataA <= 32'b00001011001110100010111011110011;
12'b000010000100: dataA <= 32'b01010000111001100011101011101000;
12'b000010000101: dataA <= 32'b00001001010111101101010000001100;
12'b000010000110: dataA <= 32'b01011010111001110110001001010011;
12'b000010000111: dataA <= 32'b00001110110111000101011000100101;
12'b000010001000: dataA <= 32'b10101101010110000011100001010000;
12'b000010001001: dataA <= 32'b00000101010110011111010001011111;
12'b000010001010: dataA <= 32'b11110000010101110010010101001010;
12'b000010001011: dataA <= 32'b00000010100101100010000100110010;
12'b000010001100: dataA <= 32'b11000101011001010110100111111000;
12'b000010001101: dataA <= 32'b00000111100101010100011011000011;
12'b000010001110: dataA <= 32'b01010001000111110010100001010001;
12'b000010001111: dataA <= 32'b00000011100011000110011111000011;
12'b000010010000: dataA <= 32'b00101000101001110011000000101011;
12'b000010010001: dataA <= 32'b00000100010000111000100000101100;
12'b000010010010: dataA <= 32'b10011011100011001110111110110111;
12'b000010010011: dataA <= 32'b00001011001101111100101010010111;
12'b000010010100: dataA <= 32'b00100100011000110011000110001001;
12'b000010010101: dataA <= 32'b00001001101010011010101100101011;
12'b000010010110: dataA <= 32'b00010011011110001110011111010011;
12'b000010010111: dataA <= 32'b00000001110100110100101101010111;
12'b000010011000: dataA <= 32'b00001001010101101110110011111010;
12'b000010011001: dataA <= 32'b00000110011110001011101001011101;
12'b000010011010: dataA <= 32'b10100000101100110110111111001110;
12'b000010011011: dataA <= 32'b00000011011011001011100001100011;
12'b000010011100: dataA <= 32'b10100101001001111010010110000001;
12'b000010011101: dataA <= 32'b00001010100011000110100101001101;
12'b000010011110: dataA <= 32'b10110011001101011111001100010111;
12'b000010011111: dataA <= 32'b00001001101000101110011000101110;
12'b000010100000: dataA <= 32'b11100111001110000001110101101000;
12'b000010100001: dataA <= 32'b00001101101111010111001111101101;
12'b000010100010: dataA <= 32'b11001101011110100010110111101101;
12'b000010100011: dataA <= 32'b00001000110001011001001111110011;
12'b000010100100: dataA <= 32'b11011111000000111111001000110101;
12'b000010100101: dataA <= 32'b00000101100111011110001010100011;
12'b000010100110: dataA <= 32'b11010011000001000101011011101111;
12'b000010100111: dataA <= 32'b00001000111011101111011101110011;
12'b000010101000: dataA <= 32'b00011000001110101100100101110100;
12'b000010101001: dataA <= 32'b00001101111001110011001010001001;
12'b000010101010: dataA <= 32'b10010111101010111111001010010101;
12'b000010101011: dataA <= 32'b00001001011110100101011010000110;
12'b000010101100: dataA <= 32'b00100111001011000101011000111000;
12'b000010101101: dataA <= 32'b00000110101000100100001000111111;
12'b000010101110: dataA <= 32'b10000010101101011100000011010010;
12'b000010101111: dataA <= 32'b00000001101000001110010100011010;
12'b000010110000: dataA <= 32'b01010010111011011110011100110010;
12'b000010110001: dataA <= 32'b00000011000100010110001101110011;
12'b000010110010: dataA <= 32'b10010101110100111100000000110000;
12'b000010110011: dataA <= 32'b00001001110011110001000010000111;
12'b000010110100: dataA <= 32'b00101010000100110100111100001001;
12'b000010110101: dataA <= 32'b00000101001101011110100010101001;
12'b000010110110: dataA <= 32'b01100001000010010101100110110111;
12'b000010110111: dataA <= 32'b00000101011101111011001001101101;
12'b000010111000: dataA <= 32'b00110110111000011011100011101011;
12'b000010111001: dataA <= 32'b00000010110111010001001111110100;
12'b000010111010: dataA <= 32'b11101110101111010101011111001111;
12'b000010111011: dataA <= 32'b00000110011110011101100010011011;
12'b000010111100: dataA <= 32'b00100000000110011111100110011101;
12'b000010111101: dataA <= 32'b00000100001010010010010000001100;
12'b000010111110: dataA <= 32'b11011011001110111100010100010111;
12'b000010111111: dataA <= 32'b00000111000010010010010001000101;
12'b000011000000: dataA <= 32'b00010100100011100110000101011010;
12'b000011000001: dataA <= 32'b00001110101000010101000000111011;
12'b000011000010: dataA <= 32'b01110000110101001100100110001110;
12'b000011000011: dataA <= 32'b00000001010001000010110001000110;
12'b000011000100: dataA <= 32'b10000100100010001001010011001010;
12'b000011000101: dataA <= 32'b00001010011110101101011101000010;
12'b000011000110: dataA <= 32'b11100010011011000111001001010110;
12'b000011000111: dataA <= 32'b00000110100001100110000101110010;
12'b000011001000: dataA <= 32'b10010111010011110101000110110010;
12'b000011001001: dataA <= 32'b00000001110100100000101110001100;
12'b000011001010: dataA <= 32'b01001111001111011110011010110111;
12'b000011001011: dataA <= 32'b00000111100100000010101110010011;
12'b000011001100: dataA <= 32'b00000111100011011100000011011010;
12'b000011001101: dataA <= 32'b00000110010110110000111010011100;
12'b000011001110: dataA <= 32'b01111010100101000011111011000010;
12'b000011001111: dataA <= 32'b00000111111000010101100101001101;
12'b000011010000: dataA <= 32'b00001100100010110101101101010010;
12'b000011010001: dataA <= 32'b00001011000110101000000101001011;
12'b000011010010: dataA <= 32'b01101110001001001110100110010110;
12'b000011010011: dataA <= 32'b00001100110001100001010010010001;
12'b000011010100: dataA <= 32'b00000101000100101011000000101110;
12'b000011010101: dataA <= 32'b00000100111101011001101001011011;
12'b000011010110: dataA <= 32'b10011111110001100100010111101101;
12'b000011010111: dataA <= 32'b00001000001000000110100001101111;
12'b000011011000: dataA <= 32'b10101100110000010100011011100011;
12'b000011011001: dataA <= 32'b00001011001101100010111011110010;
12'b000011011010: dataA <= 32'b00001110111101011011101010100111;
12'b000011011011: dataA <= 32'b00001001110111101111001000001101;
12'b000011011100: dataA <= 32'b11011010111110000110001001010011;
12'b000011011101: dataA <= 32'b00001111010100000111100000101101;
12'b000011011110: dataA <= 32'b10101111001110000011100001110011;
12'b000011011111: dataA <= 32'b00000110010111100001010001101111;
12'b000011100000: dataA <= 32'b01101010001101101010010100101011;
12'b000011100001: dataA <= 32'b00000001100111011110000100101011;
12'b000011100010: dataA <= 32'b01000111100001101110111000111000;
12'b000011100011: dataA <= 32'b00000110100101010010011110111011;
12'b000011100100: dataA <= 32'b11010001001011100010000001110100;
12'b000011100101: dataA <= 32'b00000010100101000100101010111010;
12'b000011100110: dataA <= 32'b10100110100101110011000000101110;
12'b000011100111: dataA <= 32'b00000100010001110100010100101100;
12'b000011101000: dataA <= 32'b10011101100011011110011111010100;
12'b000011101001: dataA <= 32'b00001011001100111000100010101111;
12'b000011101010: dataA <= 32'b10100000011000110011100101001010;
12'b000011101011: dataA <= 32'b00001001001010011000110000101011;
12'b000011101100: dataA <= 32'b01010111100010011110011111010000;
12'b000011101101: dataA <= 32'b00000010110111110010100101100111;
12'b000011101110: dataA <= 32'b01001011011101111110110101011100;
12'b000011101111: dataA <= 32'b00000111111110001111110001100101;
12'b000011110000: dataA <= 32'b10011110101101000111001111001011;
12'b000011110001: dataA <= 32'b00000100011101001101101001011011;
12'b000011110010: dataA <= 32'b11100111000101110010100100100010;
12'b000011110011: dataA <= 32'b00001001100010000100101101010101;
12'b000011110100: dataA <= 32'b00110011000101110111011101010101;
12'b000011110101: dataA <= 32'b00001000101000101010010100111111;
12'b000011110110: dataA <= 32'b00100111001001110001110101001001;
12'b000011110111: dataA <= 32'b00001101101101011001010011110101;
12'b000011111000: dataA <= 32'b00010001100010011010100111001101;
12'b000011111001: dataA <= 32'b00001000110001011011001111110011;
12'b000011111010: dataA <= 32'b10011111000001010111011001010101;
12'b000011111011: dataA <= 32'b00000100101001011000001110011011;
12'b000011111100: dataA <= 32'b11010101000101001101101011101110;
12'b000011111101: dataA <= 32'b00001001111010110001010101110011;
12'b000011111110: dataA <= 32'b00010010010010110100010110010101;
12'b000011111111: dataA <= 32'b00001110110110110011000001111001;
12'b000100000000: dataA <= 32'b01011101101111010110101010110100;
12'b000100000001: dataA <= 32'b00001010111110100111011010010110;
12'b000100000010: dataA <= 32'b01101001000111001100111001011000;
12'b000100000011: dataA <= 32'b00000110001000011110000101001111;
12'b000100000100: dataA <= 32'b00000010111001011100000011110100;
12'b000100000101: dataA <= 32'b00000000101010001010011100010011;
12'b000100000110: dataA <= 32'b01010011000011101101111100110000;
12'b000100000111: dataA <= 32'b00000010000110010010010001110011;
12'b000100001000: dataA <= 32'b10011011111000111100010001010011;
12'b000100001001: dataA <= 32'b00001001110011101110111010010111;
12'b000100001010: dataA <= 32'b11100100000100111101011011100111;
12'b000100001011: dataA <= 32'b00000101001110011010100010010000;
12'b000100001100: dataA <= 32'b10100001000010011101100111010111;
12'b000100001101: dataA <= 32'b00000110111110111100111101110101;
12'b000100001110: dataA <= 32'b01110110110000011100000011101100;
12'b000100001111: dataA <= 32'b00000011011001010011010111110011;
12'b000100010000: dataA <= 32'b10101100101011011100111111001101;
12'b000100010001: dataA <= 32'b00000111111110100001100010010011;
12'b000100010010: dataA <= 32'b10011010000110110111010111111101;
12'b000100010011: dataA <= 32'b00000011101100001110010100001100;
12'b000100010100: dataA <= 32'b00011101010010111100000101011000;
12'b000100010101: dataA <= 32'b00000101100010001110010101010110;
12'b000100010110: dataA <= 32'b10010010100111101101010110011010;
12'b000100010111: dataA <= 32'b00001101100110010101000100110011;
12'b000100011000: dataA <= 32'b10110000101101001100110110001110;
12'b000100011001: dataA <= 32'b00000001010100000010111101010110;
12'b000100011010: dataA <= 32'b00000010101101110001010010101100;
12'b000100011011: dataA <= 32'b00001011111101101111011000111011;
12'b000100011100: dataA <= 32'b11100000011011010110101001110110;
12'b000100011101: dataA <= 32'b00000101000001100000000101101010;
12'b000100011110: dataA <= 32'b10011001010111110100010111010010;
12'b000100011111: dataA <= 32'b00000010010110011110101110001100;
12'b000100100000: dataA <= 32'b01010001010011101101111011010110;
12'b000100100001: dataA <= 32'b00000110100101000010111010001011;
12'b000100100010: dataA <= 32'b11001011101011011011100100111100;
12'b000100100011: dataA <= 32'b00000110110110110000110110011011;
12'b000100100100: dataA <= 32'b10111000011101000100001001100001;
12'b000100100101: dataA <= 32'b00001000110111011001101001011101;
12'b000100100110: dataA <= 32'b01001010101011000101011101010000;
12'b000100100111: dataA <= 32'b00001010000101100100000101001011;
12'b000100101000: dataA <= 32'b01101000000101011110110110110110;
12'b000100101001: dataA <= 32'b00001100110000100001010010000001;
12'b000100101010: dataA <= 32'b01000101010000100011100000110001;
12'b000100101011: dataA <= 32'b00000101111110011101101101011011;
12'b000100101100: dataA <= 32'b10100101110001100100010111101101;
12'b000100101101: dataA <= 32'b00000111101000000010101010000111;
12'b000100101110: dataA <= 32'b00101010101100010101001010100001;
12'b000100101111: dataA <= 32'b00001011001100100000110111100010;
12'b000100110000: dataA <= 32'b11010001000101011011111001100110;
12'b000100110001: dataA <= 32'b00001010110110101111000100010101;
12'b000100110010: dataA <= 32'b01011010111110001110001001110010;
12'b000100110011: dataA <= 32'b00001111010001001011101000111110;
12'b000100110100: dataA <= 32'b10110001001010000011100010010101;
12'b000100110101: dataA <= 32'b00000110111000100001010010000111;
12'b000100110110: dataA <= 32'b11100110001001100010010100001101;
12'b000100110111: dataA <= 32'b00000001001010011000001000101011;
12'b000100111000: dataA <= 32'b00001011101001111111001001011000;
12'b000100111001: dataA <= 32'b00000101100110001110100010111011;
12'b000100111010: dataA <= 32'b10010011010011010001010010010110;
12'b000100111011: dataA <= 32'b00000001101000000010110110110010;
12'b000100111100: dataA <= 32'b00100100100101101011000000110001;
12'b000100111101: dataA <= 32'b00000100110010110000001100110101;
12'b000100111110: dataA <= 32'b00100001100011101101111111010001;
12'b000100111111: dataA <= 32'b00001010101011110100010110111111;
12'b000101000000: dataA <= 32'b01011100011000110100000101001011;
12'b000101000001: dataA <= 32'b00001000101001011000110000101100;
12'b000101000010: dataA <= 32'b01011001100010101110001111001101;
12'b000101000011: dataA <= 32'b00000011011001101110100001111111;
12'b000101000100: dataA <= 32'b10001111100110001110110110011101;
12'b000101000101: dataA <= 32'b00001001011110010101110101101101;
12'b000101000110: dataA <= 32'b11011110101101011111101110101000;
12'b000101000111: dataA <= 32'b00000101111110010011110001011011;
12'b000101001000: dataA <= 32'b00100111000101100010100011100011;
12'b000101001001: dataA <= 32'b00001000000010000010111001100110;
12'b000101001010: dataA <= 32'b01110010111110000111011101010011;
12'b000101001011: dataA <= 32'b00001000001000100110010001010111;
12'b000101001100: dataA <= 32'b01101001000101101001110100101011;
12'b000101001101: dataA <= 32'b00001101001011011011010011110100;
12'b000101001110: dataA <= 32'b01010101101010010010010111001101;
12'b000101001111: dataA <= 32'b00001001010000011101010011101010;
12'b000101010000: dataA <= 32'b10011111000001101111101001110100;
12'b000101010001: dataA <= 32'b00000100001010010100010010011011;
12'b000101010010: dataA <= 32'b11010101001101010110001011001101;
12'b000101010011: dataA <= 32'b00001010111001110011001101110011;
12'b000101010100: dataA <= 32'b01001110010110110011110110110110;
12'b000101010101: dataA <= 32'b00001111010011110010111001101001;
12'b000101010110: dataA <= 32'b00100001101111100110001011010011;
12'b000101010111: dataA <= 32'b00001011111100101001010110100110;
12'b000101011000: dataA <= 32'b10101001000011010100011010010111;
12'b000101011001: dataA <= 32'b00000101101001011010001001100111;
12'b000101011010: dataA <= 32'b11000011000101011100010100010110;
12'b000101011011: dataA <= 32'b00000000101101001000101000010011;
12'b000101011100: dataA <= 32'b10010011000111110101001100101111;
12'b000101011101: dataA <= 32'b00000001001000001110011001101011;
12'b000101011110: dataA <= 32'b01100001111000111100110001110110;
12'b000101011111: dataA <= 32'b00001010010010101110110110101111;
12'b000101100000: dataA <= 32'b11011110000101000101111010100110;
12'b000101100001: dataA <= 32'b00000101001111011000100110000000;
12'b000101100010: dataA <= 32'b10100001000010100101011000010111;
12'b000101100011: dataA <= 32'b00001000011110111010110101111101;
12'b000101100100: dataA <= 32'b10110100101000100100110011001110;
12'b000101100101: dataA <= 32'b00000100011010010101011011110010;
12'b000101100110: dataA <= 32'b10101010100111100100001110101010;
12'b000101100111: dataA <= 32'b00001001011110100101100010010011;
12'b000101101000: dataA <= 32'b01010110000111000111001001011101;
12'b000101101001: dataA <= 32'b00000011101110001010011100010101;
12'b000101101010: dataA <= 32'b01011111010010111011100101111001;
12'b000101101011: dataA <= 32'b00000100100011001010011101011110;
12'b000101101100: dataA <= 32'b00010000101111110100100111011011;
12'b000101101101: dataA <= 32'b00001100100100010111001000110100;
12'b000101101110: dataA <= 32'b11101110101001010101000110001111;
12'b000101101111: dataA <= 32'b00000001110110000011001001100110;
12'b000101110000: dataA <= 32'b10000010111001100001010010101110;
12'b000101110001: dataA <= 32'b00001100111011110001010000111011;
12'b000101110010: dataA <= 32'b00011100011011100101111010010101;
12'b000101110011: dataA <= 32'b00000100000011011010000101100011;
12'b000101110100: dataA <= 32'b01011011010111110011100111010010;
12'b000101110101: dataA <= 32'b00000011011000011100101110010100;
12'b000101110110: dataA <= 32'b01010011011011110101001011110100;
12'b000101110111: dataA <= 32'b00000101100101000011000110001011;
12'b000101111000: dataA <= 32'b10010001110011010011000101111101;
12'b000101111001: dataA <= 32'b00000111110111101110101110011011;
12'b000101111010: dataA <= 32'b11110100010101001100101000000001;
12'b000101111011: dataA <= 32'b00001001010111011101101001100101;
12'b000101111100: dataA <= 32'b11001000110011000100111101001110;
12'b000101111101: dataA <= 32'b00001001000101011110000101000011;
12'b000101111110: dataA <= 32'b01100010000101101111000111110111;
12'b000101111111: dataA <= 32'b00001100101110100011010001110001;
12'b000110000000: dataA <= 32'b10000111011000100100010000110100;
12'b000110000001: dataA <= 32'b00000111011110100011101101010011;
12'b000110000010: dataA <= 32'b10101001101101100100100111101101;
12'b000110000011: dataA <= 32'b00000110101001000010110110011111;
12'b000110000100: dataA <= 32'b01101000101000011101101001000001;
12'b000110000101: dataA <= 32'b00001010101011100000110111010001;
12'b000110000110: dataA <= 32'b01010001001001011100001000100101;
12'b000110000111: dataA <= 32'b00001011010101101110111100100110;
12'b000110001000: dataA <= 32'b11011011000010011110001001110001;
12'b000110001001: dataA <= 32'b00001111001110010001110001001110;
12'b000110001010: dataA <= 32'b10110001000001111011100010111000;
12'b000110001011: dataA <= 32'b00000111111000100011010010011111;
12'b000110001100: dataA <= 32'b01100000001001011010100100001110;
12'b000110001101: dataA <= 32'b00000000101101010010001100101100;
12'b000110001110: dataA <= 32'b11010001110010001110111010010111;
12'b000110001111: dataA <= 32'b00000101000111001100101010110010;
12'b000110010000: dataA <= 32'b01010101010111000000110011011000;
12'b000110010001: dataA <= 32'b00000000101010000011000010101010;
12'b000110010010: dataA <= 32'b01100000100001100011010000110100;
12'b000110010011: dataA <= 32'b00000101010100101100001000111101;
12'b000110010100: dataA <= 32'b10100101100011110101001111001110;
12'b000110010101: dataA <= 32'b00001010001010110000001111010110;
12'b000110010110: dataA <= 32'b11011000011100110100100100101101;
12'b000110010111: dataA <= 32'b00001000001001010110110100101100;
12'b000110011000: dataA <= 32'b01011101100110111101111111001010;
12'b000110011001: dataA <= 32'b00000100011010101100011010010111;
12'b000110011010: dataA <= 32'b10010011101110011110100111111101;
12'b000110011011: dataA <= 32'b00001010111110011011111001110101;
12'b000110011100: dataA <= 32'b00011100101101101111101101100110;
12'b000110011101: dataA <= 32'b00000111011110010111110101011100;
12'b000110011110: dataA <= 32'b00100111000001011010110010100101;
12'b000110011111: dataA <= 32'b00000110100010000011000101110110;
12'b000110100000: dataA <= 32'b10110010110110011111011101110001;
12'b000110100001: dataA <= 32'b00000111001000100000001101101111;
12'b000110100010: dataA <= 32'b10101001000001011010000100001100;
12'b000110100011: dataA <= 32'b00001100101001011101010111110011;
12'b000110100100: dataA <= 32'b11011001101110001010010110101110;
12'b000110100101: dataA <= 32'b00001001010000011111010011100001;
12'b000110100110: dataA <= 32'b01011111000010000111101010010011;
12'b000110100111: dataA <= 32'b00000011101011001110010110011011;
12'b000110101000: dataA <= 32'b00010111010001100110001010101011;
12'b000110101001: dataA <= 32'b00001011111000110101000101110100;
12'b000110101010: dataA <= 32'b01001010011110110011100111010110;
12'b000110101011: dataA <= 32'b00001111010000110000110001011001;
12'b000110101100: dataA <= 32'b11100101101111101101101011110010;
12'b000110101101: dataA <= 32'b00001101011010101011010010110101;
12'b000110101110: dataA <= 32'b10101001000011010011111010110110;
12'b000110101111: dataA <= 32'b00000100101010010100001001111111;
12'b000110110000: dataA <= 32'b01000011010001100100100100110111;
12'b000110110001: dataA <= 32'b00000000110000000110110000010100;
12'b000110110010: dataA <= 32'b10010101001011110100011100101101;
12'b000110110011: dataA <= 32'b00000000101011001010100001101011;
12'b000110110100: dataA <= 32'b00100111111001000101010010011000;
12'b000110110101: dataA <= 32'b00001010010001101100101111000111;
12'b000110110110: dataA <= 32'b11011000000101010110001001100101;
12'b000110110111: dataA <= 32'b00000101010000010110101001101000;
12'b000110111000: dataA <= 32'b10100001000010101101001000110111;
12'b000110111001: dataA <= 32'b00001001111110111010101010001101;
12'b000110111010: dataA <= 32'b00110000100000101101010011010000;
12'b000110111011: dataA <= 32'b00000101011011011001011111100010;
12'b000110111100: dataA <= 32'b01101000100011100011101110000111;
12'b000110111101: dataA <= 32'b00001010011110100111011110010011;
12'b000110111110: dataA <= 32'b00010000001111010110101010011100;
12'b000110111111: dataA <= 32'b00000011101111001000100100011110;
12'b000111000000: dataA <= 32'b10011111010010111011010110111010;
12'b000111000001: dataA <= 32'b00000011000101001000100101101110;
12'b000111000010: dataA <= 32'b01001110110011110100001000011011;
12'b000111000011: dataA <= 32'b00001011100010010111001100110100;
12'b000111000100: dataA <= 32'b00101100100101011101010110010000;
12'b000111000101: dataA <= 32'b00000010111001000101010101111111;
12'b000111000110: dataA <= 32'b11000011000101010001100010110001;
12'b000111000111: dataA <= 32'b00001101111001110011001000111011;
12'b000111001000: dataA <= 32'b00011000011111110101011010110100;
12'b000111001001: dataA <= 32'b00000010100101010100001001100011;
12'b000111001010: dataA <= 32'b01011101011011110010110111110011;
12'b000111001011: dataA <= 32'b00000100011010011010101110010100;
12'b000111001100: dataA <= 32'b00010101011111110100011100010011;
12'b000111001101: dataA <= 32'b00000100100110000011010010000011;
12'b000111001110: dataA <= 32'b10010101111011010010100111011101;
12'b000111001111: dataA <= 32'b00001000010111101100101010011011;
12'b000111010000: dataA <= 32'b11101110001101001100110110100001;
12'b000111010001: dataA <= 32'b00001010010110100011101001101101;
12'b000111010010: dataA <= 32'b00000110111111001100011100101100;
12'b000111010011: dataA <= 32'b00001000000100011000000101000100;
12'b000111010100: dataA <= 32'b10011100000110000111001000010111;
12'b000111010101: dataA <= 32'b00001100001100100101001101100001;
12'b000111010110: dataA <= 32'b11001011100100101100110001010110;
12'b000111010111: dataA <= 32'b00001000111110100111101001010011;
12'b000111011000: dataA <= 32'b01101101101001101100110111001110;
12'b000111011001: dataA <= 32'b00000110001001000011000010110111;
12'b000111011010: dataA <= 32'b11100110100100101110010111100001;
12'b000111011011: dataA <= 32'b00001010001010100000110111000000;
12'b000111011100: dataA <= 32'b11010011010001011100010111100101;
12'b000111011101: dataA <= 32'b00001011110011101110111000110110;
12'b000111011110: dataA <= 32'b00011011000010101101111001110001;
12'b000111011111: dataA <= 32'b00001111001011010101111001011111;
12'b000111100000: dataA <= 32'b01110000111001111011100011111010;
12'b000111100001: dataA <= 32'b00001000111000100101001110110111;
12'b000111100010: dataA <= 32'b11011100001001010010110011110000;
12'b000111100011: dataA <= 32'b00000000101111001110010000110100;
12'b000111100100: dataA <= 32'b01010101111010100110111010110110;
12'b000111100101: dataA <= 32'b00000100001000001010110010101010;
12'b000111100110: dataA <= 32'b00010111011010110000100100011010;
12'b000111100111: dataA <= 32'b00000000101101000011001110100010;
12'b000111101000: dataA <= 32'b11011110100001100011100001010110;
12'b000111101001: dataA <= 32'b00000101010101100110000101000101;
12'b000111101010: dataA <= 32'b00100111011111110100011111001011;
12'b000111101011: dataA <= 32'b00001001101001101100001011100110;
12'b000111101100: dataA <= 32'b01010110011100110101000100001110;
12'b000111101101: dataA <= 32'b00000111001001010110111000110101;
12'b000111101110: dataA <= 32'b00100001100111000101011110001000;
12'b000111101111: dataA <= 32'b00000101011011101000010110100111;
12'b000111110000: dataA <= 32'b10010111110010101110101000111101;
12'b000111110001: dataA <= 32'b00001011111100100001111001111101;
12'b000111110010: dataA <= 32'b01011010110010000111101100100100;
12'b000111110011: dataA <= 32'b00001000111110011101110101011100;
12'b000111110100: dataA <= 32'b00100110111101011011000001101000;
12'b000111110101: dataA <= 32'b00000101100011000101010001111110;
12'b000111110110: dataA <= 32'b10110010101110101111001101101111;
12'b000111110111: dataA <= 32'b00000110101000011100001101111111;
12'b000111111000: dataA <= 32'b11101001000001010010010100001101;
12'b000111111001: dataA <= 32'b00001011100111011111010111110010;
12'b000111111010: dataA <= 32'b01011101101110000010010110101110;
12'b000111111011: dataA <= 32'b00001001010000011111010011010001;
12'b000111111100: dataA <= 32'b00011111000010011111101010110010;
12'b000111111101: dataA <= 32'b00000011101101001010011110010011;
12'b000111111110: dataA <= 32'b00011001010001110110011010101010;
12'b000111111111: dataA <= 32'b00001100010110110100111101110100;
12'b001000000000: dataA <= 32'b10001000100110101011010111110110;
12'b001000000001: dataA <= 32'b00001111001101110000101101001001;
12'b001000000010: dataA <= 32'b10101001101011110100111011110000;
12'b001000000011: dataA <= 32'b00001110011000101101001110111101;
12'b001000000100: dataA <= 32'b10101000111111010011011011010101;
12'b001000000101: dataA <= 32'b00000100001011010000010010010111;
12'b001000000110: dataA <= 32'b00000101011101100100110101111000;
12'b001000000111: dataA <= 32'b00000000110011000100111100011101;
12'b001000001000: dataA <= 32'b11010101001111110011101100001011;
12'b001000001001: dataA <= 32'b00000000101110001000101001101011;
12'b001000001010: dataA <= 32'b10101011110101001101100011011010;
12'b001000001011: dataA <= 32'b00001010110000101010101011010110;
12'b001000001100: dataA <= 32'b00010010001001100110011000100100;
12'b001000001101: dataA <= 32'b00000101010001010100101101011001;
12'b001000001110: dataA <= 32'b01100001000010110100101001110111;
12'b001000001111: dataA <= 32'b00001010111101110110100010010101;
12'b001000010000: dataA <= 32'b01101110011000110101110011010010;
12'b001000010001: dataA <= 32'b00000110111100011011011111011001;
12'b001000010010: dataA <= 32'b01100100011111011011001101000101;
12'b001000010011: dataA <= 32'b00001011111100101011011010001011;
12'b001000010100: dataA <= 32'b10001100010011100101111011011011;
12'b001000010101: dataA <= 32'b00000011110001000110110000101110;
12'b001000010110: dataA <= 32'b10100001010010110010110111111010;
12'b001000010111: dataA <= 32'b00000010100111000110110001111110;
12'b001000011000: dataA <= 32'b11001110111011110011011001011011;
12'b001000011001: dataA <= 32'b00001010000001011001010000111100;
12'b001000011010: dataA <= 32'b11101000011101101101100110010001;
12'b001000011011: dataA <= 32'b00000011111010000111100010001110;
12'b001000011100: dataA <= 32'b01000011010001001001110010110011;
12'b001000011101: dataA <= 32'b00001110110111110101000000111100;
12'b001000011110: dataA <= 32'b01010110100011110100101011010010;
12'b001000011111: dataA <= 32'b00000001100111001110001101011011;
12'b001000100000: dataA <= 32'b00100001011011101010001000010011;
12'b001000100001: dataA <= 32'b00000101011011011010101110010100;
12'b001000100010: dataA <= 32'b00011001100011110011101100010001;
12'b001000100011: dataA <= 32'b00000011101000000101011101111011;
12'b001000100100: dataA <= 32'b01011011111011000010001000111101;
12'b001000100101: dataA <= 32'b00001001010110101010100110010011;
12'b001000100110: dataA <= 32'b00101010000101010101000101100001;
12'b001000100111: dataA <= 32'b00001010110101100111101001111110;
12'b001000101000: dataA <= 32'b10001001000111001011111100101010;
12'b001000101001: dataA <= 32'b00000111000100010010001001001100;
12'b001000101010: dataA <= 32'b10010110000110010111001001010110;
12'b001000101011: dataA <= 32'b00001011101011100111001101010001;
12'b001000101100: dataA <= 32'b00001111101000110101010010011001;
12'b001000101101: dataA <= 32'b00001010011110101011100101010100;
12'b001000101110: dataA <= 32'b11110001100001101100110111001110;
12'b001000101111: dataA <= 32'b00000101101010000011001111001110;
12'b001000110000: dataA <= 32'b10100100100100111110100110000001;
12'b001000110001: dataA <= 32'b00001001001001011110110110110000;
12'b001000110010: dataA <= 32'b01010101010101100100010110100101;
12'b001000110011: dataA <= 32'b00001011110010101110110001000111;
12'b001000110100: dataA <= 32'b01011011000110110101101010010000;
12'b001000110101: dataA <= 32'b00001110101000011011111001110111;
12'b001000110110: dataA <= 32'b11110000110101111011100100111011;
12'b001000110111: dataA <= 32'b00001001011000100111001111001110;
12'b001000111000: dataA <= 32'b01010110001101001011010100010001;
12'b001000111001: dataA <= 32'b00000000110010001010011000110101;
12'b001000111010: dataA <= 32'b00011011111010110110101011010101;
12'b001000111011: dataA <= 32'b00000011101010001000111010100010;
12'b001000111100: dataA <= 32'b11011001011110011000010101011011;
12'b001000111101: dataA <= 32'b00000000110000000101010110010001;
12'b001000111110: dataA <= 32'b00011010100101100011100010011001;
12'b001000111111: dataA <= 32'b00000110010110100000000101010110;
12'b001001000000: dataA <= 32'b10101011011011110011101110101000;
12'b001001000001: dataA <= 32'b00001001001001100110000111101101;
12'b001001000010: dataA <= 32'b10010010100000111101010100001111;
12'b001001000011: dataA <= 32'b00000110101010010100111100111101;
12'b001001000100: dataA <= 32'b11100101100111001100111101100101;
12'b001001000101: dataA <= 32'b00000110111100100100010110110110;
12'b001001000110: dataA <= 32'b10011101110110111110001010011100;
12'b001001000111: dataA <= 32'b00001101011011100101111010001101;
12'b001001001000: dataA <= 32'b01011000110010011111101011100010;
12'b001001001001: dataA <= 32'b00001010011110100011110101100100;
12'b001001001010: dataA <= 32'b00100110111001010011010000101010;
12'b001001001011: dataA <= 32'b00000100100100000111011010001110;
12'b001001001100: dataA <= 32'b10110000101011000110101101101101;
12'b001001001101: dataA <= 32'b00000101101001011000010010010111;
12'b001001001110: dataA <= 32'b00101000111101001010100011101111;
12'b001001001111: dataA <= 32'b00001011000110100001010111101010;
12'b001001010000: dataA <= 32'b11100001101101110010010110101111;
12'b001001010001: dataA <= 32'b00001001001111100001010010111000;
12'b001001010010: dataA <= 32'b00011111000010101111011010110001;
12'b001001010011: dataA <= 32'b00000011001111001000100110010011;
12'b001001010100: dataA <= 32'b00011011010110000110011001101001;
12'b001001010101: dataA <= 32'b00001100110101110100110101110100;
12'b001001010110: dataA <= 32'b00000110110010101011001000110110;
12'b001001010111: dataA <= 32'b00001111001011101110100100111010;
12'b001001011000: dataA <= 32'b00101101100111110100001011101111;
12'b001001011001: dataA <= 32'b00001110110110101101001011000101;
12'b001001011010: dataA <= 32'b10101000111011001010111011110011;
12'b001001011011: dataA <= 32'b00000100001101001010010110100111;
12'b001001011100: dataA <= 32'b10001001100101101100110110111001;
12'b001001011101: dataA <= 32'b00000001010110000101000100100101;
12'b001001011110: dataA <= 32'b11010111010011110010111011101001;
12'b001001011111: dataA <= 32'b00000000110001000110110001101011;
12'b001001100000: dataA <= 32'b00110001110001011101110100011100;
12'b001001100001: dataA <= 32'b00001010101111101000100111100110;
12'b001001100010: dataA <= 32'b01001110001101110110010111100100;
12'b001001100011: dataA <= 32'b00000101010010010010110001001001;
12'b001001100100: dataA <= 32'b01100001000010110100011010010110;
12'b001001100101: dataA <= 32'b00001100011100110100010110011101;
12'b001001100110: dataA <= 32'b11101010010101000110010011110100;
12'b001001100111: dataA <= 32'b00000111111101011111011111000000;
12'b001001101000: dataA <= 32'b01100000011111010010101100000011;
12'b001001101001: dataA <= 32'b00001100111011101101010110001011;
12'b001001101010: dataA <= 32'b00001000011011110101011100111001;
12'b001001101011: dataA <= 32'b00000011110011000110111000111111;
12'b001001101100: dataA <= 32'b10100011010010101010101001011010;
12'b001001101101: dataA <= 32'b00000001101001000110111010010110;
12'b001001101110: dataA <= 32'b01001101000011101010101010011010;
12'b001001101111: dataA <= 32'b00001000100001011011010001000101;
12'b001001110000: dataA <= 32'b11100100011101110101100110010001;
12'b001001110001: dataA <= 32'b00000100111100001011101010011110;
12'b001001110010: dataA <= 32'b11000101011100111010010011010101;
12'b001001110011: dataA <= 32'b00001111010100110100111000111100;
12'b001001110100: dataA <= 32'b10010010100111110011111011010001;
12'b001001110101: dataA <= 32'b00000001001001001010010101011011;
12'b001001110110: dataA <= 32'b00100011011011011001101000010011;
12'b001001110111: dataA <= 32'b00000110011100011000110010010100;
12'b001001111000: dataA <= 32'b00011101100011110010111100101111;
12'b001001111001: dataA <= 32'b00000011001010001001100101111011;
12'b001001111010: dataA <= 32'b01100001111010110001101001111101;
12'b001001111011: dataA <= 32'b00001001110110100110100010010011;
12'b001001111100: dataA <= 32'b00100100000101011101010100000011;
12'b001001111101: dataA <= 32'b00001011010100101011100110001110;
12'b001001111110: dataA <= 32'b11001001001111001011011011101000;
12'b001001111111: dataA <= 32'b00000110000101001110010001001100;
12'b001010000000: dataA <= 32'b00010000001010100110111001110110;
12'b001010000001: dataA <= 32'b00001011001001100111001001000010;
12'b001010000010: dataA <= 32'b01010011110000111101110011011011;
12'b001010000011: dataA <= 32'b00001011111101101111100001010100;
12'b001010000100: dataA <= 32'b10110101011101110100110111001110;
12'b001010000101: dataA <= 32'b00000101001011000101011011011110;
12'b001010000110: dataA <= 32'b01100000100101001111000100100010;
12'b001010000111: dataA <= 32'b00001000101001011110110110011000;
12'b001010001000: dataA <= 32'b10010111011001100100100101100110;
12'b001010001001: dataA <= 32'b00001011110000101100101101011111;
12'b001010001010: dataA <= 32'b01011011000110111101001010001111;
12'b001010001011: dataA <= 32'b00001101100110100001111010000111;
12'b001010001100: dataA <= 32'b10101110101101111011100101111100;
12'b001010001101: dataA <= 32'b00001010010111100111001011011110;
12'b001010001110: dataA <= 32'b11010010010001001011100100010011;
12'b001010001111: dataA <= 32'b00000001010101000110100001000101;
12'b001010010000: dataA <= 32'b00100001111011000110001011110011;
12'b001010010001: dataA <= 32'b00000011001100001001000010010010;
12'b001010010010: dataA <= 32'b11011101011110000000010110011100;
12'b001010010011: dataA <= 32'b00000000110011000111100010000001;
12'b001010010100: dataA <= 32'b01011000100101100011110011011011;
12'b001010010101: dataA <= 32'b00000110110110011010000101100110;
12'b001010010110: dataA <= 32'b11101101010111110010111101100110;
12'b001010010111: dataA <= 32'b00001000001001100000000111110100;
12'b001010011000: dataA <= 32'b00010000101001001101110100010001;
12'b001010011001: dataA <= 32'b00000110001010010101000001001110;
12'b001010011010: dataA <= 32'b01101001100011001100011100000011;
12'b001010011011: dataA <= 32'b00000111111101100000010011001110;
12'b001010011100: dataA <= 32'b10100001110111001101101011011011;
12'b001010011101: dataA <= 32'b00001110011000101011110110010101;
12'b001010011110: dataA <= 32'b10011000110110110111011010000001;
12'b001010011111: dataA <= 32'b00001011111101100111110101100100;
12'b001010100000: dataA <= 32'b00100110111001010011100000101101;
12'b001010100001: dataA <= 32'b00000011000110001011100010011110;
12'b001010100010: dataA <= 32'b01101100100011010110011101001011;
12'b001010100011: dataA <= 32'b00000101001010010100010110101111;
12'b001010100100: dataA <= 32'b10101000111001000011000011110001;
12'b001010100101: dataA <= 32'b00001010000101100011010111011001;
12'b001010100110: dataA <= 32'b01100101101101101010010110101111;
12'b001010100111: dataA <= 32'b00001001001111100011010010101000;
12'b001010101000: dataA <= 32'b00011111000011000111001010110000;
12'b001010101001: dataA <= 32'b00000011010001000110101110001011;
12'b001010101010: dataA <= 32'b00011101010110010110011001001001;
12'b001010101011: dataA <= 32'b00001101010011110010101101110100;
12'b001010101100: dataA <= 32'b10000110111010100010111001010110;
12'b001010101101: dataA <= 32'b00001110001000101010100000110010;
12'b001010101110: dataA <= 32'b10110001011111110011011011101101;
12'b001010101111: dataA <= 32'b00001111010011101101000011001100;
12'b001010110000: dataA <= 32'b11011100101101011001101001101000;
12'b001010110001: dataA <= 32'b00000110110111001011101011110010;
12'b001010110010: dataA <= 32'b11110011101110011100101100110010;
12'b001010110011: dataA <= 32'b00001011011101100011110110110110;
12'b001010110100: dataA <= 32'b10101001010001011000010100101000;
12'b001010110101: dataA <= 32'b00001000111110011001110001111100;
12'b001010110110: dataA <= 32'b11111000011110111101001110010111;
12'b001010110111: dataA <= 32'b00000111101010010010101111000000;
12'b001010111000: dataA <= 32'b10000111100011001100010010010000;
12'b001010111001: dataA <= 32'b00001001010101011001011000101101;
12'b001010111010: dataA <= 32'b00100000111110001010011011001011;
12'b001010111011: dataA <= 32'b00001110000111001010010110101011;
12'b001010111100: dataA <= 32'b11001010101011001101111010011000;
12'b001010111101: dataA <= 32'b00001110110000101111000000011001;
12'b001010111110: dataA <= 32'b10001110111101010001010001100111;
12'b001010111111: dataA <= 32'b00001101100110101010100101101011;
12'b001011000000: dataA <= 32'b00001101101110101000011100100110;
12'b001011000001: dataA <= 32'b00001001111000011101110011100110;
12'b001011000010: dataA <= 32'b01101000111001010010101101001101;
12'b001011000011: dataA <= 32'b00000100111100011101110011010011;
12'b001011000100: dataA <= 32'b11100001100101010000101101001011;
12'b001011000101: dataA <= 32'b00000000101110101001001010101101;
12'b001011000110: dataA <= 32'b00001110110110110100011000110011;
12'b001011000111: dataA <= 32'b00001110010110110101101011011011;
12'b001011001000: dataA <= 32'b00101111110101001110001010111001;
12'b001011001001: dataA <= 32'b00001010000001011100010110011110;
12'b001011001010: dataA <= 32'b00010011011001111000011000101001;
12'b001011001011: dataA <= 32'b00000100111101001011101001110101;
12'b001011001100: dataA <= 32'b01101100111000110001001001101111;
12'b001011001101: dataA <= 32'b00001110010011011001001110000011;
12'b001011001110: dataA <= 32'b00110001000101011000010111100110;
12'b001011001111: dataA <= 32'b00000101011001110011101101100100;
12'b001011010000: dataA <= 32'b01111100111100110010011110101100;
12'b001011010001: dataA <= 32'b00001011001100010000110001101011;
12'b001011010010: dataA <= 32'b10000010110110101101000001110111;
12'b001011010011: dataA <= 32'b00001010001001110010101011000011;
12'b001011010100: dataA <= 32'b10100111101101101001100100001000;
12'b001011010101: dataA <= 32'b00000010110011001001100010011101;
12'b001011010110: dataA <= 32'b11000101011111011010111011001100;
12'b001011010111: dataA <= 32'b00000100101001100100110001000101;
12'b001011011000: dataA <= 32'b01111001011010111110001101111001;
12'b001011011001: dataA <= 32'b00001110101000110000100010001101;
12'b001011011010: dataA <= 32'b00101110010110011100010111010001;
12'b001011011011: dataA <= 32'b00000101110101101101110111010001;
12'b001011011100: dataA <= 32'b00010010111111100101100001010110;
12'b001011011101: dataA <= 32'b00000100101110011011000000001011;
12'b001011011110: dataA <= 32'b00101101010010010100110011010100;
12'b001011011111: dataA <= 32'b00001000001000010110100111110101;
12'b001011100000: dataA <= 32'b11100011001010100010000111101011;
12'b001011100001: dataA <= 32'b00000011000100111100111111101011;
12'b001011100010: dataA <= 32'b00010110100001110100001110010100;
12'b001011100011: dataA <= 32'b00001011101011100100110011010001;
12'b001011100100: dataA <= 32'b11001001011001110101101001110111;
12'b001011100101: dataA <= 32'b00001010111101010001110010111101;
12'b001011100110: dataA <= 32'b01111100111111000001111001101000;
12'b001011100111: dataA <= 32'b00000110011001100001101101000011;
12'b001011101000: dataA <= 32'b11101111000100001011111110010011;
12'b001011101001: dataA <= 32'b00001001111110110001110000111011;
12'b001011101010: dataA <= 32'b11010011001101111100111101111001;
12'b001011101011: dataA <= 32'b00001011010010000011001011001100;
12'b001011101100: dataA <= 32'b01101010100101011000010011000100;
12'b001011101101: dataA <= 32'b00000100101111000010111110011000;
12'b001011101110: dataA <= 32'b10010101011110111101101000110111;
12'b001011101111: dataA <= 32'b00000101010011100001010111000101;
12'b001011110000: dataA <= 32'b10110000101110001001100001100111;
12'b001011110001: dataA <= 32'b00001110110000001000111111001001;
12'b001011110010: dataA <= 32'b01111010111110110001101101101001;
12'b001011110011: dataA <= 32'b00001100000011111010101010110011;
12'b001011110100: dataA <= 32'b11011011001111101010010000101011;
12'b001011110101: dataA <= 32'b00001110101000111010110010010100;
12'b001011110110: dataA <= 32'b00011100110001110101010110111110;
12'b001011110111: dataA <= 32'b00000011011001110001101011000011;
12'b001011111000: dataA <= 32'b10010000100111001001010101100101;
12'b001011111001: dataA <= 32'b00000101010101001011010111101010;
12'b001011111010: dataA <= 32'b00011100101101100101111000111000;
12'b001011111011: dataA <= 32'b00000010101011101010111000110001;
12'b001011111100: dataA <= 32'b10110110110101001100100111110010;
12'b001011111101: dataA <= 32'b00000111101101101000111000001010;
12'b001011111110: dataA <= 32'b10100001000011100001111000001010;
12'b001011111111: dataA <= 32'b00001000111001010111110001100011;
12'b001100000000: dataA <= 32'b01101011000111001011010100101101;
12'b001100000001: dataA <= 32'b00001001100101010110011010000100;
12'b001100000010: dataA <= 32'b01011101110001011010111011001101;
12'b001100000011: dataA <= 32'b00000100000011010000101001010110;
12'b001100000100: dataA <= 32'b10101110011101101000010110101000;
12'b001100000101: dataA <= 32'b00001001100001100000100110010001;
12'b001100000110: dataA <= 32'b01011110101101101001011010101001;
12'b001100000111: dataA <= 32'b00000101110111001001011111110011;
12'b001100001000: dataA <= 32'b00101111110110011100111100010100;
12'b001100001001: dataA <= 32'b00001001111110011111110110100111;
12'b001100001010: dataA <= 32'b10100111010101110000010101100111;
12'b001100001011: dataA <= 32'b00000111011110010101101101111100;
12'b001100001100: dataA <= 32'b01111010101010110101101101011001;
12'b001100001101: dataA <= 32'b00001000001010010100101011010001;
12'b001100001110: dataA <= 32'b00000101011011001100110010001110;
12'b001100001111: dataA <= 32'b00001000110101010111010100100101;
12'b001100010000: dataA <= 32'b01100000111110010010011011101100;
12'b001100010001: dataA <= 32'b00001110101010010000010010101011;
12'b001100010010: dataA <= 32'b00001100100010111110011001011001;
12'b001100010011: dataA <= 32'b00001110010010101111001000101001;
12'b001100010100: dataA <= 32'b10001110110101100001000010100101;
12'b001100010101: dataA <= 32'b00001110001000101100101001101011;
12'b001100010110: dataA <= 32'b10001001100110111000111101101001;
12'b001100010111: dataA <= 32'b00001000111000011001110011010110;
12'b001100011000: dataA <= 32'b00101000111101011010011101010000;
12'b001100011001: dataA <= 32'b00000011111010011001110011010100;
12'b001100011010: dataA <= 32'b00011101100001101000011101101101;
12'b001100011011: dataA <= 32'b00000000101011101001001110011110;
12'b001100011100: dataA <= 32'b10001110101110110100101000110011;
12'b001100011101: dataA <= 32'b00001101011000110001110011011011;
12'b001100011110: dataA <= 32'b00101001111000111101101001111010;
12'b001100011111: dataA <= 32'b00001011100010100000010110001110;
12'b001100100000: dataA <= 32'b00010001010010010000011001001001;
12'b001100100001: dataA <= 32'b00000011111100000111100001101101;
12'b001100100010: dataA <= 32'b01101100111101000000101001101111;
12'b001100100011: dataA <= 32'b00001101110101010111001010000011;
12'b001100100100: dataA <= 32'b00110001001101110000011000100111;
12'b001100100101: dataA <= 32'b00000100011000101111110101100100;
12'b001100100110: dataA <= 32'b01111101001001000001111110101110;
12'b001100100111: dataA <= 32'b00001011001101010010101001101011;
12'b001100101000: dataA <= 32'b00000010101010100101010000110100;
12'b001100101001: dataA <= 32'b00001010101010110100110011000100;
12'b001100101010: dataA <= 32'b10100011101101111001100101000110;
12'b001100101011: dataA <= 32'b00000010010001000101011010010101;
12'b001100101100: dataA <= 32'b01000011010011100011011011001101;
12'b001100101101: dataA <= 32'b00000101101000100110110000110101;
12'b001100101110: dataA <= 32'b01110101100010101110011100111011;
12'b001100101111: dataA <= 32'b00001111001011110010101010000101;
12'b001100110000: dataA <= 32'b10110000011110011100100111010001;
12'b001100110001: dataA <= 32'b00000101010100100111111011011001;
12'b001100110010: dataA <= 32'b01010010110111010110000000110011;
12'b001100110011: dataA <= 32'b00000100101101011011000000010010;
12'b001100110100: dataA <= 32'b11101011010110001100110010110010;
12'b001100110101: dataA <= 32'b00001001001000011000100011101101;
12'b001100110110: dataA <= 32'b01100011001010110010011000001011;
12'b001100110111: dataA <= 32'b00000100000010111101001011101100;
12'b001100111000: dataA <= 32'b10011010011101110100001101110110;
12'b001100111001: dataA <= 32'b00001100001101100110110011011001;
12'b001100111010: dataA <= 32'b01000111010001101101101000110111;
12'b001100111011: dataA <= 32'b00001001011110001101101010101110;
12'b001100111100: dataA <= 32'b11111101001011010010011010101001;
12'b001100111101: dataA <= 32'b00000101011000011101101101000010;
12'b001100111110: dataA <= 32'b01101111001100001011001101110101;
12'b001100111111: dataA <= 32'b00001000011110101011110100111011;
12'b001101000000: dataA <= 32'b01010011001001110100111100111011;
12'b001101000001: dataA <= 32'b00001011010011000010111111000101;
12'b001101000010: dataA <= 32'b10101100101001110000010100000010;
12'b001101000011: dataA <= 32'b00000100101101000010110010110000;
12'b001101000100: dataA <= 32'b00010001011010101110000111110111;
12'b001101000101: dataA <= 32'b00000101010010011111010110110110;
12'b001101000110: dataA <= 32'b01110010110110011001100010100100;
12'b001101000111: dataA <= 32'b00001110010010001010110111011010;
12'b001101001000: dataA <= 32'b10111011000111000010001110001011;
12'b001101001001: dataA <= 32'b00001101100101111100110110110011;
12'b001101001010: dataA <= 32'b11011001001111110011000001001000;
12'b001101001011: dataA <= 32'b00001111001011111010111010001100;
12'b001101001100: dataA <= 32'b10011100110001101101010101011110;
12'b001101001101: dataA <= 32'b00000010010110101101110011000011;
12'b001101001110: dataA <= 32'b01010100011111010001110110100100;
12'b001101001111: dataA <= 32'b00000100110100001001001111110011;
12'b001101010000: dataA <= 32'b10011110101101010101100111111000;
12'b001101010001: dataA <= 32'b00000011001001101010111101000000;
12'b001101010010: dataA <= 32'b00110110111101001100010111110010;
12'b001101010011: dataA <= 32'b00000111101101101000111100011010;
12'b001101010100: dataA <= 32'b01100001000011101010101000101010;
12'b001101010101: dataA <= 32'b00000111111001010011101101100011;
12'b001101010110: dataA <= 32'b01101011001011001011110100101100;
12'b001101010111: dataA <= 32'b00001010100110011010010110000100;
12'b001101011000: dataA <= 32'b00011001110001100010101011001110;
12'b001101011001: dataA <= 32'b00000101100001010010100001000110;
12'b001101011010: dataA <= 32'b11110010100110000000010111101000;
12'b001101011011: dataA <= 32'b00001011000010100100100110100001;
12'b001101011100: dataA <= 32'b00100000101101111001011011001010;
12'b001101011101: dataA <= 32'b00000101010110000101010111110100;
12'b001101011110: dataA <= 32'b01101001111010010100111011110110;
12'b001101011111: dataA <= 32'b00001000011110011001110010001111;
12'b001101100000: dataA <= 32'b10100101010110001000010110100110;
12'b001101100001: dataA <= 32'b00000101111110010001101001110100;
12'b001101100010: dataA <= 32'b11111100110010101101111100011011;
12'b001101100011: dataA <= 32'b00001000101011010110100111100001;
12'b001101100100: dataA <= 32'b10000011001111000101010010101100;
12'b001101100101: dataA <= 32'b00001000010101010101010000011100;
12'b001101100110: dataA <= 32'b10100000111110100010101011101110;
12'b001101100111: dataA <= 32'b00001111001100010100001010110011;
12'b001101101000: dataA <= 32'b11010000011110101110101000011001;
12'b001101101001: dataA <= 32'b00001101110101101111001101000000;
12'b001101101010: dataA <= 32'b01010000101101110000110011100011;
12'b001101101011: dataA <= 32'b00001111001011101110110001101011;
12'b001101101100: dataA <= 32'b00000111011111010001011110001011;
12'b001101101101: dataA <= 32'b00000111111000010011101111000111;
12'b001101101110: dataA <= 32'b10101001000001101010001101010010;
12'b001101101111: dataA <= 32'b00000010111001010011101111010100;
12'b001101110000: dataA <= 32'b01011001100010000000011101101111;
12'b001101110001: dataA <= 32'b00000001001000100111010010001110;
12'b001101110010: dataA <= 32'b00010010100110101101001000010011;
12'b001101110011: dataA <= 32'b00001100111010101011110111100100;
12'b001101110100: dataA <= 32'b00100011111000110101011000111010;
12'b001101110101: dataA <= 32'b00001100100100100100011001111110;
12'b001101110110: dataA <= 32'b11001111001110101000011010001010;
12'b001101110111: dataA <= 32'b00000010111010000101010101100100;
12'b001101111000: dataA <= 32'b01101101000101011000011001110000;
12'b001101111001: dataA <= 32'b00001101010111010111001010001011;
12'b001101111010: dataA <= 32'b11101111010110001000011001100111;
12'b001101111011: dataA <= 32'b00000011010110101001111001100011;
12'b001101111100: dataA <= 32'b00111101010101010001011110110001;
12'b001101111101: dataA <= 32'b00001011101111010100100101110011;
12'b001101111110: dataA <= 32'b10000110100010011101100000110010;
12'b001101111111: dataA <= 32'b00001011001011110100111010111100;
12'b001110000000: dataA <= 32'b11011111110010001001100110000110;
12'b001110000001: dataA <= 32'b00000010001111000011001110000101;
12'b001110000010: dataA <= 32'b11000011000111100011111011101111;
12'b001110000011: dataA <= 32'b00000110000111100110110100110100;
12'b001110000100: dataA <= 32'b01110011101010011110101011011101;
12'b001110000101: dataA <= 32'b00001111001110110100110001111101;
12'b001110000110: dataA <= 32'b01110100100110011100100111010001;
12'b001110000111: dataA <= 32'b00000100110011100001111011101010;
12'b001110001000: dataA <= 32'b11010010110011001110100000110000;
12'b001110001001: dataA <= 32'b00000101001011011010111100011001;
12'b001110001010: dataA <= 32'b01101001011010001101000010110000;
12'b001110001011: dataA <= 32'b00001001101000011100100011011110;
12'b001110001100: dataA <= 32'b00100001001010111010101000101100;
12'b001110001101: dataA <= 32'b00000101100001111101010111100101;
12'b001110001110: dataA <= 32'b01011100011101110100001101011000;
12'b001110001111: dataA <= 32'b00001100001110100110110111101010;
12'b001110010000: dataA <= 32'b01000101000101011101011000011000;
12'b001110010001: dataA <= 32'b00000111111110001001100010011110;
12'b001110010010: dataA <= 32'b10111101010111011010111011001010;
12'b001110010011: dataA <= 32'b00000100010111011001101001001010;
12'b001110010100: dataA <= 32'b11101101010000010010011101010111;
12'b001110010101: dataA <= 32'b00000110111110100111111001000010;
12'b001110010110: dataA <= 32'b11010001000001110100111011011101;
12'b001110010111: dataA <= 32'b00001010110101000010110010111101;
12'b001110011000: dataA <= 32'b11101110110010001000010101100001;
12'b001110011001: dataA <= 32'b00000100101100000100100111000000;
12'b001110011010: dataA <= 32'b01001111010010100110010111010111;
12'b001110011011: dataA <= 32'b00000100110001011101010010101110;
12'b001110011100: dataA <= 32'b11110010111110101001110100000011;
12'b001110011101: dataA <= 32'b00001101110101001010101111100010;
12'b001110011110: dataA <= 32'b00111001010011010010101110101110;
12'b001110011111: dataA <= 32'b00001110001000111100111110110100;
12'b001110100000: dataA <= 32'b00011001001011110011110010000110;
12'b001110100001: dataA <= 32'b00001111001110111011000110001101;
12'b001110100010: dataA <= 32'b00011110110001100101000100011100;
12'b001110100011: dataA <= 32'b00000001110100101001110111000100;
12'b001110100100: dataA <= 32'b00010110011011100010100111100100;
12'b001110100101: dataA <= 32'b00000100010010000111000111110100;
12'b001110100110: dataA <= 32'b01100000101101001101010110110111;
12'b001110100111: dataA <= 32'b00000011101000101011000001011000;
12'b001110101000: dataA <= 32'b01110111000101001011110111010010;
12'b001110101001: dataA <= 32'b00001000001101101001000000101001;
12'b001110101010: dataA <= 32'b01100001000011110011001001001010;
12'b001110101011: dataA <= 32'b00000110111000001111101001100011;
12'b001110101100: dataA <= 32'b01101001001111001100010101001010;
12'b001110101101: dataA <= 32'b00001011000111011110010110000100;
12'b001110101110: dataA <= 32'b10010011101101101010101011010000;
12'b001110101111: dataA <= 32'b00000110100001010110011100110101;
12'b001110110000: dataA <= 32'b00110100101110011000011000001000;
12'b001110110001: dataA <= 32'b00001100000011100110100110110010;
12'b001110110010: dataA <= 32'b11100000101110001001011011101011;
12'b001110110011: dataA <= 32'b00000100110100000101001011110100;
12'b001110110100: dataA <= 32'b01100011111010001101001011010111;
12'b001110110101: dataA <= 32'b00000110111110010101101101111111;
12'b001110110110: dataA <= 32'b10100011011010100000010111100110;
12'b001110110111: dataA <= 32'b00000100011101001101100001110100;
12'b001110111000: dataA <= 32'b10111100111110011110001011011100;
12'b001110111001: dataA <= 32'b00001001001011011010100011101010;
12'b001110111010: dataA <= 32'b11000011000010111101110011001010;
12'b001110111011: dataA <= 32'b00000111110101010011001100011011;
12'b001110111100: dataA <= 32'b00100000111110101010111011101111;
12'b001110111101: dataA <= 32'b00001111001111011010001010110100;
12'b001110111110: dataA <= 32'b01010100010110011110110111011001;
12'b001110111111: dataA <= 32'b00001101010111101101010101010000;
12'b001111000000: dataA <= 32'b01010010101010000000110101000010;
12'b001111000001: dataA <= 32'b00001111001101110000110101110011;
12'b001111000010: dataA <= 32'b01000011010011100001111110101101;
12'b001111000011: dataA <= 32'b00000111011000001111101010101111;
12'b001111000100: dataA <= 32'b00101001000001110010001100110100;
12'b001111000101: dataA <= 32'b00000001110110001111101011001101;
12'b001111000110: dataA <= 32'b01010111011110010000011101110001;
12'b001111000111: dataA <= 32'b00000010000110100101010010000110;
12'b001111001000: dataA <= 32'b11010100100010100101010111110011;
12'b001111001001: dataA <= 32'b00001011011100100101111011011100;
12'b001111001010: dataA <= 32'b00011101111000101100110111011010;
12'b001111001011: dataA <= 32'b00001101100110101000011101110110;
12'b001111001100: dataA <= 32'b11001101000110111000111010101011;
12'b001111001101: dataA <= 32'b00000001110111000011001001100100;
12'b001111001110: dataA <= 32'b01101011001001110000011001010001;
12'b001111001111: dataA <= 32'b00001100011001010111000110001011;
12'b001111010000: dataA <= 32'b10101101011010100000011010001000;
12'b001111010001: dataA <= 32'b00000010110100100011111001101011;
12'b001111010010: dataA <= 32'b00111001011101100001011110110100;
12'b001111010011: dataA <= 32'b00001011110000010110100001110011;
12'b001111010100: dataA <= 32'b11001010010110010101100000101111;
12'b001111010101: dataA <= 32'b00001011101101110101000110111100;
12'b001111010110: dataA <= 32'b11011001101110011001110111000101;
12'b001111010111: dataA <= 32'b00000010101101000011000001111101;
12'b001111011000: dataA <= 32'b01000010111011100100101011110000;
12'b001111011001: dataA <= 32'b00000111000110101000111000101100;
12'b001111011010: dataA <= 32'b01101101110010001110111010011110;
12'b001111011011: dataA <= 32'b00001111010001110110111001110101;
12'b001111011100: dataA <= 32'b00110110101110010100110110110000;
12'b001111011101: dataA <= 32'b00000100110010011011111011110011;
12'b001111011110: dataA <= 32'b01010100101110110111000000101101;
12'b001111011111: dataA <= 32'b00000101101010011010111100101001;
12'b001111100000: dataA <= 32'b11100101011110000101000010101110;
12'b001111100001: dataA <= 32'b00001010101001011110100011001110;
12'b001111100010: dataA <= 32'b10100001001011000011001000101100;
12'b001111100011: dataA <= 32'b00000111000001111001011111011101;
12'b001111100100: dataA <= 32'b00100000011101110100001100011010;
12'b001111100101: dataA <= 32'b00001100010000101000111011110011;
12'b001111100110: dataA <= 32'b10000100111101010101000111010111;
12'b001111100111: dataA <= 32'b00000110111110000111011010001110;
12'b001111101000: dataA <= 32'b01111001011111011011101011101011;
12'b001111101001: dataA <= 32'b00000011110101010101100101011010;
12'b001111101010: dataA <= 32'b10101011010100011001111100011001;
12'b001111101011: dataA <= 32'b00000101011110100001111001001010;
12'b001111101100: dataA <= 32'b00010000111101101100111010011110;
12'b001111101101: dataA <= 32'b00001010010101000100100110101110;
12'b001111101110: dataA <= 32'b01110000110110100000010111000001;
12'b001111101111: dataA <= 32'b00000101001011000110011111010001;
12'b001111110000: dataA <= 32'b10001111001110010110010110110110;
12'b001111110001: dataA <= 32'b00000100101111011011010010011110;
12'b001111110010: dataA <= 32'b01110011000110111010000101000001;
12'b001111110011: dataA <= 32'b00001101010111001100100111101011;
12'b001111110100: dataA <= 32'b01110111011011010011001110110000;
12'b001111110101: dataA <= 32'b00001111001010111101001010110100;
12'b001111110110: dataA <= 32'b00010111000111110100100011000100;
12'b001111110111: dataA <= 32'b00001111010001111011010010000101;
12'b001111111000: dataA <= 32'b01100000110001011101000010111010;
12'b001111111001: dataA <= 32'b00000001010010100011111011000100;
12'b001111111010: dataA <= 32'b10011010011011101011001000100100;
12'b001111111011: dataA <= 32'b00000100010001000110111111110100;
12'b001111111100: dataA <= 32'b01100000101101000101000110010111;
12'b001111111101: dataA <= 32'b00000100100110101011000101110000;
12'b001111111110: dataA <= 32'b11110111001101001011100111010010;
12'b001111111111: dataA <= 32'b00001000001101101001000000111000;
12'b010000000000: dataA <= 32'b00100001000011110011111001101011;
12'b010000000001: dataA <= 32'b00000101111000001011100001101011;
12'b010000000010: dataA <= 32'b01101001010011000100110101101010;
12'b010000000011: dataA <= 32'b00001100001000100010010110000100;
12'b010000000100: dataA <= 32'b00001111101001110010011011010001;
12'b010000000101: dataA <= 32'b00001000000001011000011100101101;
12'b010000000110: dataA <= 32'b01110110110110110000101001001000;
12'b010000000111: dataA <= 32'b00001101000101101000101010111010;
12'b010000001000: dataA <= 32'b10100010101110011001101100001101;
12'b010000001001: dataA <= 32'b00000100010011000011000011101101;
12'b010000001010: dataA <= 32'b01011101111010000101001010011000;
12'b010000001011: dataA <= 32'b00000101011110001111101001100111;
12'b010000001100: dataA <= 32'b01100001011010111000101000000110;
12'b010000001101: dataA <= 32'b00000011011011001001011001101100;
12'b010000001110: dataA <= 32'b01111101001010001110001001111101;
12'b010000001111: dataA <= 32'b00001001101100011100100011110011;
12'b010000010000: dataA <= 32'b01000010110110101110000011101000;
12'b010000010001: dataA <= 32'b00000111010101010001001000011011;
12'b010000010010: dataA <= 32'b01100000111110110011001011110001;
12'b010000010011: dataA <= 32'b00001111010010011110000110110100;
12'b010000010100: dataA <= 32'b01011000010010000111000110011000;
12'b010000010101: dataA <= 32'b00001100111001101011011001101000;
12'b010000010110: dataA <= 32'b01010100100110011001000110100001;
12'b010000010111: dataA <= 32'b00001111010000110000111101110011;
12'b010000011000: dataA <= 32'b10000011001011101010011110110000;
12'b010000011001: dataA <= 32'b00000110011000001011100010010111;
12'b010000011010: dataA <= 32'b01101001000110000010001100010101;
12'b010000011011: dataA <= 32'b00000001010100001011100011000101;
12'b010000011100: dataA <= 32'b01010011011010101000101101010011;
12'b010000011101: dataA <= 32'b00000011000100100011010101110110;
12'b010000011110: dataA <= 32'b01010110011110011101100111010011;
12'b010000011111: dataA <= 32'b00001010011101011111111011010101;
12'b010000100000: dataA <= 32'b00010111111000101100010110011010;
12'b010000100001: dataA <= 32'b00001110101000101100100001100110;
12'b010000100010: dataA <= 32'b10001100111111010001011011001100;
12'b010000100011: dataA <= 32'b00000000110101000010111101011100;
12'b010000100100: dataA <= 32'b10101011001110001000011001010001;
12'b010000100101: dataA <= 32'b00001011011011010111000010010011;
12'b010000100110: dataA <= 32'b10101001011110111000101011001001;
12'b010000100111: dataA <= 32'b00000010110010011101111001101011;
12'b010000101000: dataA <= 32'b00110101101001110001001110010110;
12'b010000101001: dataA <= 32'b00001011010010011010011101111011;
12'b010000101010: dataA <= 32'b00001110001110000101110000101100;
12'b010000101011: dataA <= 32'b00001011101110110101001110110101;
12'b010000101100: dataA <= 32'b10010101101010101001111000000101;
12'b010000101101: dataA <= 32'b00000010101011000010110101101101;
12'b010000101110: dataA <= 32'b11000010101111011101001011010010;
12'b010000101111: dataA <= 32'b00001000000110101000111100101011;
12'b010000110000: dataA <= 32'b00101001110101110110111000111110;
12'b010000110001: dataA <= 32'b00001111010100110111000101101101;
12'b010000110010: dataA <= 32'b11111000110110001100110110110000;
12'b010000110011: dataA <= 32'b00000100010000010101111011110011;
12'b010000110100: dataA <= 32'b11010110101010100111010000101010;
12'b010000110101: dataA <= 32'b00000110001001011010111101000000;
12'b010000110110: dataA <= 32'b01100011011101111101000011001100;
12'b010000110111: dataA <= 32'b00001011001010100010100010111111;
12'b010000111000: dataA <= 32'b00011111001011000011101001001100;
12'b010000111001: dataA <= 32'b00001000100001110101101011001110;
12'b010000111010: dataA <= 32'b11100100011101110011111010111011;
12'b010000111011: dataA <= 32'b00001100010010101000111111110011;
12'b010000111100: dataA <= 32'b10000100110001001100110110110111;
12'b010000111101: dataA <= 32'b00000101011101000101001101111110;
12'b010000111110: dataA <= 32'b00110101101011100100001100001101;
12'b010000111111: dataA <= 32'b00000011010100010001100001100010;
12'b010001000000: dataA <= 32'b01101001011000101001011011011011;
12'b010001000001: dataA <= 32'b00000100011100011011111001010010;
12'b010001000010: dataA <= 32'b01010010110101100100101000111110;
12'b010001000011: dataA <= 32'b00001001010110000110011110100110;
12'b010001000100: dataA <= 32'b00110000111110111000101000100001;
12'b010001000101: dataA <= 32'b00000101101010001010010111100010;
12'b010001000110: dataA <= 32'b10001101000110000110010101110101;
12'b010001000111: dataA <= 32'b00000100101110011001001110001110;
12'b010001001000: dataA <= 32'b00110001001111000010100110100001;
12'b010001001001: dataA <= 32'b00001100111001010000100011101100;
12'b010001001010: dataA <= 32'b10110011100011011011101110110011;
12'b010001001011: dataA <= 32'b00001111001101111011010110110100;
12'b010001001100: dataA <= 32'b00010111000011110101000100000010;
12'b010001001101: dataA <= 32'b00001111010100111001011001111101;
12'b010001001110: dataA <= 32'b11100010110001010100110001111000;
12'b010001001111: dataA <= 32'b00000001001111011101111011000100;
12'b010001010000: dataA <= 32'b01011110011011101011111001100101;
12'b010001010001: dataA <= 32'b00000100001111001000110011101101;
12'b010001010010: dataA <= 32'b01100010101100111100100101110110;
12'b010001010011: dataA <= 32'b00000101100101101001001010001000;
12'b010001010100: dataA <= 32'b10110101010101001011010110110001;
12'b010001010101: dataA <= 32'b00001000001101101001000101001000;
12'b010001010110: dataA <= 32'b00100001000011110100101010001100;
12'b010001010111: dataA <= 32'b00000101010111001001010101110011;
12'b010001011000: dataA <= 32'b01100111010111000101010110101001;
12'b010001011001: dataA <= 32'b00001100101010100110011001111100;
12'b010001011010: dataA <= 32'b10001011100001111010011011010010;
12'b010001011011: dataA <= 32'b00001001100001011100011000101100;
12'b010001011100: dataA <= 32'b11110110111111000000111001101001;
12'b010001011101: dataA <= 32'b00001110001000101010101111000010;
12'b010001011110: dataA <= 32'b00100100110010101001111100001110;
12'b010001011111: dataA <= 32'b00000100010010000100110111100110;
12'b010001100000: dataA <= 32'b00010111111010000101001001011001;
12'b010001100001: dataA <= 32'b00000100011100001011100001010111;
12'b010001100010: dataA <= 32'b01011101011011001001001001000110;
12'b010001100011: dataA <= 32'b00000010011001000111010001101100;
12'b010001100100: dataA <= 32'b11111011010110000110001000011110;
12'b010001100101: dataA <= 32'b00001001101100100000011111110011;
12'b010001100110: dataA <= 32'b10000010101010011110010100100111;
12'b010001100111: dataA <= 32'b00000110110101010001000000100010;
12'b010001101000: dataA <= 32'b10100000111110110011011011110010;
12'b010001101001: dataA <= 32'b00001110110101100100001010101100;
12'b010001101010: dataA <= 32'b01011100010001110111000101111000;
12'b010001101011: dataA <= 32'b00001011111010100111011110000000;
12'b010001101100: dataA <= 32'b00010110100010101001010111100001;
12'b010001101101: dataA <= 32'b00001111010011110001000101111011;
12'b010001101110: dataA <= 32'b10000010111111110011001110110011;
12'b010001101111: dataA <= 32'b00000101010111001001011010000111;
12'b010001110000: dataA <= 32'b11100111001010001010001011110111;
12'b010001110001: dataA <= 32'b00000001010001001001011010111101;
12'b010001110010: dataA <= 32'b00010001010111000000111101010101;
12'b010001110011: dataA <= 32'b00000100000010100001010101100110;
12'b010001110100: dataA <= 32'b11011010011110010101100111010011;
12'b010001110101: dataA <= 32'b00001000111101011001111011001101;
12'b010001110110: dataA <= 32'b11010001110100101011100101011001;
12'b010001110111: dataA <= 32'b00001111001011101110100101010101;
12'b010001111000: dataA <= 32'b01001100111011100001111011001101;
12'b010001111001: dataA <= 32'b00000000110010000010110001011100;
12'b010001111010: dataA <= 32'b10101001010010100000011001010010;
12'b010001111011: dataA <= 32'b00001010011100010110111110010011;
12'b010001111100: dataA <= 32'b01100111100011001001001011101010;
12'b010001111101: dataA <= 32'b00000010010000010111111001101011;
12'b010001111110: dataA <= 32'b00110001110010000001001101011001;
12'b010001111111: dataA <= 32'b00001011010011011100011110000011;
12'b010010000000: dataA <= 32'b10010010001001111101110001001001;
12'b010010000001: dataA <= 32'b00001100010000110011010110101101;
12'b010010000010: dataA <= 32'b10010001100110110010011001000101;
12'b010010000011: dataA <= 32'b00000011001001000010101101100101;
12'b010010000100: dataA <= 32'b01000100100011010101101011010011;
12'b010010000101: dataA <= 32'b00001000100110101000111100101011;
12'b010010000110: dataA <= 32'b00100011110101100110100111011110;
12'b010010000111: dataA <= 32'b00001110110110110101001101100101;
12'b010010001000: dataA <= 32'b10111001000010001100110110110000;
12'b010010001001: dataA <= 32'b00000100001111010001110011110100;
12'b010010001010: dataA <= 32'b01011000100110001111010001101000;
12'b010010001011: dataA <= 32'b00000110101001011100111001010000;
12'b010010001100: dataA <= 32'b10011111100001110101000011101010;
12'b010010001101: dataA <= 32'b00001011101100100100100010100111;
12'b010010001110: dataA <= 32'b10011111001011000011111001101101;
12'b010010001111: dataA <= 32'b00001010000001110001110010111110;
12'b010010010000: dataA <= 32'b10100110100001110011111001111100;
12'b010010010001: dataA <= 32'b00001011110011101000111111110100;
12'b010010010010: dataA <= 32'b10000110101001001100100101110110;
12'b010010010011: dataA <= 32'b00000011111100000011000001101110;
12'b010010010100: dataA <= 32'b00110001110011011100101100001110;
12'b010010010101: dataA <= 32'b00000010110010001111011001101010;
12'b010010010110: dataA <= 32'b00100101011101000000111010011100;
12'b010010010111: dataA <= 32'b00000010111010010101110101011010;
12'b010010011000: dataA <= 32'b10010010110001100100010111011110;
12'b010010011001: dataA <= 32'b00001000110111001010010110010110;
12'b010010011010: dataA <= 32'b10110001000111001001001010000001;
12'b010010011011: dataA <= 32'b00000110001001010000001111110010;
12'b010010011100: dataA <= 32'b10001100111101110110010101010101;
12'b010010011101: dataA <= 32'b00000101001101011001001101110110;
12'b010010011110: dataA <= 32'b11110001010011001011001000000001;
12'b010010011111: dataA <= 32'b00001011111010010010011011101100;
12'b010010100000: dataA <= 32'b11101111101011011100001110010101;
12'b010010100001: dataA <= 32'b00001111010000111001100010101100;
12'b010010100010: dataA <= 32'b00010111000011100101110101100001;
12'b010010100011: dataA <= 32'b00001110110111110101100101110101;
12'b010010100100: dataA <= 32'b01100010110001010100010001010110;
12'b010010100101: dataA <= 32'b00000001001100010111110110111101;
12'b010010100110: dataA <= 32'b00100010011011101100011010100101;
12'b010010100111: dataA <= 32'b00000100001110001010101011100110;
12'b010010101000: dataA <= 32'b01100100110000111100010100110101;
12'b010010101001: dataA <= 32'b00000110100100101001001110100000;
12'b010010101010: dataA <= 32'b01110001011101010011000110110001;
12'b010010101011: dataA <= 32'b00001000101110100111001001100000;
12'b010010101100: dataA <= 32'b00100001000011101101011010101101;
12'b010010101101: dataA <= 32'b00000100110110000111001101110011;
12'b010010101110: dataA <= 32'b01100011010110110101100111001000;
12'b010010101111: dataA <= 32'b00001101001100101010011101111100;
12'b010010110000: dataA <= 32'b00001001011010001010011010110011;
12'b010010110001: dataA <= 32'b00001011000010100000011000100100;
12'b010010110010: dataA <= 32'b01110111000111010001011010001010;
12'b010010110011: dataA <= 32'b00001111001010101100110011001011;
12'b010010110100: dataA <= 32'b11100110110010111010001100010000;
12'b010010110101: dataA <= 32'b00000011110000000100101011010110;
12'b010010110110: dataA <= 32'b10010001110101111101001000011010;
12'b010010110111: dataA <= 32'b00000010111011001001011000111110;
12'b010010111000: dataA <= 32'b00011011010111011001101010000111;
12'b010010111001: dataA <= 32'b00000001010111000101000101101100;
12'b010010111010: dataA <= 32'b10111001100001110110000111011110;
12'b010010111011: dataA <= 32'b00001010001101100010100011110100;
12'b010010111100: dataA <= 32'b00000110100010001110010101000110;
12'b010010111101: dataA <= 32'b00000110010100010000111100101010;
12'b010010111110: dataA <= 32'b11100000111110110011101011010100;
12'b010010111111: dataA <= 32'b00001110011000101010001010101100;
12'b010011000000: dataA <= 32'b01100000010001100110110100110111;
12'b010011000001: dataA <= 32'b00001010011100100101011110011000;
12'b010011000010: dataA <= 32'b00011010011110111001101001000001;
12'b010011000011: dataA <= 32'b00001110110110110001001010000011;
12'b010011000100: dataA <= 32'b10000010110011110011111110010101;
12'b010011000101: dataA <= 32'b00000100110110000111001101101111;
12'b010011000110: dataA <= 32'b00100111001110011010001010111000;
12'b010011000111: dataA <= 32'b00000001001110000111001110101110;
12'b010011001000: dataA <= 32'b11001111001111010001011100010111;
12'b010011001001: dataA <= 32'b00000101100001011111010101011101;
12'b010011001010: dataA <= 32'b01011110011010001101100110110010;
12'b010011001011: dataA <= 32'b00000111011101010101110110111110;
12'b010011001100: dataA <= 32'b10001101101100101011000100111000;
12'b010011001101: dataA <= 32'b00001111001110110000101101001101;
12'b010011001110: dataA <= 32'b00001110110011101010011011001110;
12'b010011001111: dataA <= 32'b00000000101111000100101001010100;
12'b010011010000: dataA <= 32'b11100111010110111000101000110010;
12'b010011010001: dataA <= 32'b00001000111101010110111010010011;
12'b010011010010: dataA <= 32'b01100011100011011001101100001100;
12'b010011010011: dataA <= 32'b00000010001110010001110101110011;
12'b010011010100: dataA <= 32'b00101101110110010001001100011010;
12'b010011010101: dataA <= 32'b00001010110100100000011110001011;
12'b010011010110: dataA <= 32'b11011000000101101101100010000110;
12'b010011010111: dataA <= 32'b00001011110001110001011010100101;
12'b010011011000: dataA <= 32'b01001101011110111010101010000110;
12'b010011011001: dataA <= 32'b00000100000111000110100001011101;
12'b010011011010: dataA <= 32'b11001000011011000110001010110100;
12'b010011011011: dataA <= 32'b00001001100111101001000000110010;
12'b010011011100: dataA <= 32'b11011101110101010110010101111110;
12'b010011011101: dataA <= 32'b00001101111001110011010101011100;
12'b010011011110: dataA <= 32'b00111001001010000101000110101111;
12'b010011011111: dataA <= 32'b00000100101101001011101111110101;
12'b010011100000: dataA <= 32'b01011010100101110111010010000101;
12'b010011100001: dataA <= 32'b00000111001001011100111001101000;
12'b010011100010: dataA <= 32'b10011101011101110100110100001000;
12'b010011100011: dataA <= 32'b00001011101101101000100110001111;
12'b010011100100: dataA <= 32'b11011101001011000100011001101101;
12'b010011100101: dataA <= 32'b00001011100010101101110110101110;
12'b010011100110: dataA <= 32'b00101010100101110011111000011101;
12'b010011100111: dataA <= 32'b00001011010101101001000011110101;
12'b010011101000: dataA <= 32'b01001010011101001100010101010101;
12'b010011101001: dataA <= 32'b00000010111010000010111001011110;
12'b010011101010: dataA <= 32'b11101101110111010101011100010000;
12'b010011101011: dataA <= 32'b00000010110000001101010101111001;
12'b010011101100: dataA <= 32'b11100011011101010000011000111101;
12'b010011101101: dataA <= 32'b00000001111000001111110001101001;
12'b010011101110: dataA <= 32'b10010100101101100100010101111110;
12'b010011101111: dataA <= 32'b00001000010111010000001110000110;
12'b010011110000: dataA <= 32'b01110001001011011001101011100010;
12'b010011110001: dataA <= 32'b00000110101001010100000111110011;
12'b010011110010: dataA <= 32'b10001100110101100110010100110011;
12'b010011110011: dataA <= 32'b00000101001100010111001001100110;
12'b010011110100: dataA <= 32'b01101111011011001011101001100001;
12'b010011110101: dataA <= 32'b00001010011100010110010111100101;
12'b010011110110: dataA <= 32'b00101011101111011100101101011000;
12'b010011110111: dataA <= 32'b00001111010011110101101010100101;
12'b010011111000: dataA <= 32'b11010110111111011110010111000001;
12'b010011111001: dataA <= 32'b00001101111001110001101001110100;
12'b010011111010: dataA <= 32'b10100100110101001100000000110011;
12'b010011111011: dataA <= 32'b00000001101010010011110010110101;
12'b010011111100: dataA <= 32'b10100110011011100101001011100111;
12'b010011111101: dataA <= 32'b00000100001100001100100011010110;
12'b010011111110: dataA <= 32'b10100110110000111011110100010100;
12'b010011111111: dataA <= 32'b00000111100100100111010010111000;
12'b010100000000: dataA <= 32'b01101111100101011010110110110000;
12'b010100000001: dataA <= 32'b00001000101110100111001101111000;
12'b010100000010: dataA <= 32'b11100001000011100110001010101110;
12'b010100000011: dataA <= 32'b00000011110100000101000001111010;
12'b010100000100: dataA <= 32'b01100001011010101101110111101000;
12'b010100000101: dataA <= 32'b00001101101110101110100001111100;
12'b010100000110: dataA <= 32'b10000111001110010010101010010100;
12'b010100000111: dataA <= 32'b00001100100100100100011000100011;
12'b010100001000: dataA <= 32'b11110101010011100010001010101011;
12'b010100001001: dataA <= 32'b00001111001101101100110111010011;
12'b010100001010: dataA <= 32'b00100110110111000010101100010010;
12'b010100001011: dataA <= 32'b00000011101110001000100010111111;
12'b010100001100: dataA <= 32'b01001101101101110101000111011010;
12'b010100001101: dataA <= 32'b00000001111000000111010000101110;
12'b010100001110: dataA <= 32'b00011001010111101010011011001000;
12'b010100001111: dataA <= 32'b00000000110100000100111101101100;
12'b010100010000: dataA <= 32'b01110101101001100110000101111101;
12'b010100010001: dataA <= 32'b00001010001110100110100011101101;
12'b010100010010: dataA <= 32'b10001010010101111110100110000101;
12'b010100010011: dataA <= 32'b00000101110011010000110100111001;
12'b010100010100: dataA <= 32'b00100000111110111100001010110101;
12'b010100010101: dataA <= 32'b00001101011010101110010010100101;
12'b010100010110: dataA <= 32'b10100100010001010110100100010101;
12'b010100010111: dataA <= 32'b00001001011100100001011110110000;
12'b010100011000: dataA <= 32'b00011110011111001010001010100010;
12'b010100011001: dataA <= 32'b00001101111000101111010010000011;
12'b010100011010: dataA <= 32'b01000100100111110100101101010111;
12'b010100011011: dataA <= 32'b00000100010100000111000101010111;
12'b010100011100: dataA <= 32'b01100101001110100010011001111001;
12'b010100011101: dataA <= 32'b00000001001100000111000110011110;
12'b010100011110: dataA <= 32'b10001111000111100001111011011001;
12'b010100011111: dataA <= 32'b00000111000001011101010101001101;
12'b010100100000: dataA <= 32'b10100010011001111101110110110010;
12'b010100100001: dataA <= 32'b00000110011101001111110010110110;
12'b010100100010: dataA <= 32'b00001001100100110010100011110110;
12'b010100100011: dataA <= 32'b00001111010001110010110101000101;
12'b010100100100: dataA <= 32'b11010000101011110011001011110000;
12'b010100100101: dataA <= 32'b00000000101100000110011101010011;
12'b010100100110: dataA <= 32'b11100101010111001001001000110010;
12'b010100100111: dataA <= 32'b00000111111101010110110110010011;
12'b010100101000: dataA <= 32'b01011111100111101010011100001110;
12'b010100101001: dataA <= 32'b00000010101100001101101101110011;
12'b010100101010: dataA <= 32'b00100111111010100001011011011100;
12'b010100101011: dataA <= 32'b00001010010101100100011110001011;
12'b010100101100: dataA <= 32'b11011110000101100101100010100100;
12'b010100101101: dataA <= 32'b00001011110011101101100010010101;
12'b010100101110: dataA <= 32'b00001011011011000011001011000111;
12'b010100101111: dataA <= 32'b00000101000110001000011001010101;
12'b010100110000: dataA <= 32'b01001100010010111110101010010101;
12'b010100110001: dataA <= 32'b00001010101000101001000100111010;
12'b010100110010: dataA <= 32'b10011001110101000110000100011101;
12'b010100110011: dataA <= 32'b00001100111011110001011101011100;
12'b010100110100: dataA <= 32'b11110111010001111101000110101111;
12'b010100110101: dataA <= 32'b00000100101100000111100011100101;
12'b010100110110: dataA <= 32'b01011110100101100111010011100011;
12'b010100110111: dataA <= 32'b00001000001000011100111010000000;
12'b010100111000: dataA <= 32'b10011001011101101100110101000111;
12'b010100111001: dataA <= 32'b00001011101111101010101001110111;
12'b010100111010: dataA <= 32'b00011101001011000100111001101110;
12'b010100111011: dataA <= 32'b00001100100100100111111010011111;
12'b010100111100: dataA <= 32'b11101100101001110011110111011101;
12'b010100111101: dataA <= 32'b00001010110110101001000111100101;
12'b010100111110: dataA <= 32'b00001100010101000011110100110100;
12'b010100111111: dataA <= 32'b00000001111000000100101101001110;
12'b010101000000: dataA <= 32'b11100111111011001101111100010010;
12'b010101000001: dataA <= 32'b00000010101101001011001110001001;
12'b010101000010: dataA <= 32'b11011111100001101000010111111101;
12'b010101000011: dataA <= 32'b00000001010110001011101001111001;
12'b010101000100: dataA <= 32'b10010110101001100100000100011101;
12'b010101000101: dataA <= 32'b00000111010111010100000101101110;
12'b010101000110: dataA <= 32'b00101111010011101010011100100100;
12'b010101000111: dataA <= 32'b00000111101001011010000111110100;
12'b010101001000: dataA <= 32'b01001110101101010110000100110010;
12'b010101001001: dataA <= 32'b00000101101011010111000101010110;
12'b010101001010: dataA <= 32'b11101011011111010100001011000010;
12'b010101001011: dataA <= 32'b00001001011100011010010111010101;
12'b010101001100: dataA <= 32'b01100111110011010101001100111010;
12'b010101001101: dataA <= 32'b00001110110110110001110010011101;
12'b010101001110: dataA <= 32'b11010110111011001110111000100001;
12'b010101001111: dataA <= 32'b00001100111011101101110001101100;
12'b010101010000: dataA <= 32'b11100100110101001011110000110000;
12'b010101010001: dataA <= 32'b00000010101000001111101010100101;
12'b010101010010: dataA <= 32'b00101010011111011101101100101001;
12'b010101010011: dataA <= 32'b00000100101011010000011011000111;
12'b010101010100: dataA <= 32'b00100110110100111011010100010010;
12'b010101010101: dataA <= 32'b00001000100100100101010011001001;
12'b010101010110: dataA <= 32'b01101011101001100010100110110000;
12'b010101010111: dataA <= 32'b00001000101110100101001110010000;
12'b010101011000: dataA <= 32'b11100001000011010110101010101111;
12'b010101011001: dataA <= 32'b00000011110010000100111010000010;
12'b010101011010: dataA <= 32'b01011111011010011110001000101000;
12'b010101011011: dataA <= 32'b00001101110000110000101001111100;
12'b010101011100: dataA <= 32'b00000111000110011010101001110101;
12'b010101011101: dataA <= 32'b00001101100101101000011100101011;
12'b010101011110: dataA <= 32'b01110011011011110010101011001100;
12'b010101011111: dataA <= 32'b00001111010000101100111111010100;
12'b010101100000: dataA <= 32'b00011010110001010001111001000111;
12'b010101100001: dataA <= 32'b00000111011000010001101111100010;
12'b010101100010: dataA <= 32'b10110111100110100100011101010001;
12'b010101100011: dataA <= 32'b00001100011100101001110011001110;
12'b010101100100: dataA <= 32'b10101011001101001000100100001001;
12'b010101100101: dataA <= 32'b00001010011110011111110110000100;
12'b010101100110: dataA <= 32'b10110100010111000100111110110100;
12'b010101100111: dataA <= 32'b00000111001011010000110010101000;
12'b010101101000: dataA <= 32'b00001011101011010100000010110011;
12'b010101101001: dataA <= 32'b00001001110100011011011100110110;
12'b010101101010: dataA <= 32'b11011110111110000010001010101010;
12'b010101101011: dataA <= 32'b00001101000101001000100010100010;
12'b010101101100: dataA <= 32'b01001000110111010101011010110111;
12'b010101101101: dataA <= 32'b00001110001101101110111100010010;
12'b010101101110: dataA <= 32'b11001111000001000001100001001010;
12'b010101101111: dataA <= 32'b00001100000100101000100001100011;
12'b010101110000: dataA <= 32'b01010011110110010000011011100101;
12'b010101110001: dataA <= 32'b00001010010111100011110011101101;
12'b010101110010: dataA <= 32'b00100110110101001010111100101100;
12'b010101110011: dataA <= 32'b00000110011101100011110011001011;
12'b010101110100: dataA <= 32'b10100011100000111000111100101001;
12'b010101110101: dataA <= 32'b00000000110001101011000110110101;
12'b010101110110: dataA <= 32'b01001100111010111100001001010010;
12'b010101110111: dataA <= 32'b00001110110011111001100011010010;
12'b010101111000: dataA <= 32'b11110011101101010110011011011000;
12'b010101111001: dataA <= 32'b00001000100001011010011010100101;
12'b010101111010: dataA <= 32'b01010101011101100000011000001000;
12'b010101111011: dataA <= 32'b00000110011110001111110001111101;
12'b010101111100: dataA <= 32'b01101010110100100001101001001110;
12'b010101111101: dataA <= 32'b00001110110000011011010001111011;
12'b010101111110: dataA <= 32'b01110011000001001000100111000111;
12'b010101111111: dataA <= 32'b00000110011010110111100101101100;
12'b010110000000: dataA <= 32'b10111100110000101010111110001001;
12'b010110000001: dataA <= 32'b00001010101011001110110101100011;
12'b010110000010: dataA <= 32'b01000011000010110100110010011010;
12'b010110000011: dataA <= 32'b00001001101000110000100110111011;
12'b010110000100: dataA <= 32'b01101101101001100001110011101001;
12'b010110000101: dataA <= 32'b00000011010101001101101110100101;
12'b010110000110: dataA <= 32'b00001001100111010010001010101011;
12'b010110000111: dataA <= 32'b00000100001010100010101101001110;
12'b010110001000: dataA <= 32'b00111011001111000101111110110111;
12'b010110001001: dataA <= 32'b00001101100110101110011110010101;
12'b010110001010: dataA <= 32'b11101000010010100100000111110010;
12'b010110001011: dataA <= 32'b00000110010110110001110010111000;
12'b010110001100: dataA <= 32'b11010011000011101100110001111000;
12'b010110001101: dataA <= 32'b00000100001111011101000100001011;
12'b010110001110: dataA <= 32'b01101111001110011100100011110101;
12'b010110001111: dataA <= 32'b00000111101000010100101011110100;
12'b010110010000: dataA <= 32'b00100101000110011001110111001100;
12'b010110010001: dataA <= 32'b00000010000110111100110011100011;
12'b010110010010: dataA <= 32'b11010100100101111100011110110001;
12'b010110010011: dataA <= 32'b00001011001010100010101110111000;
12'b010110010100: dataA <= 32'b10001011100101111101111010010110;
12'b010110010101: dataA <= 32'b00001100011100010111110111000101;
12'b010110010110: dataA <= 32'b10111100110010111001101001000111;
12'b010110010111: dataA <= 32'b00000110111010100111101000111011;
12'b010110011000: dataA <= 32'b00110001000000001100101110110000;
12'b010110011001: dataA <= 32'b00001011011101110101101000111100;
12'b010110011010: dataA <= 32'b10010101010010000100111110110111;
12'b010110011011: dataA <= 32'b00001011110001000011010111010100;
12'b010110011100: dataA <= 32'b01101000100001001000100010000110;
12'b010110011101: dataA <= 32'b00000100110000000011001010000000;
12'b010110011110: dataA <= 32'b01010111100011000101011001010110;
12'b010110011111: dataA <= 32'b00000101110100100011010011001101;
12'b010110100000: dataA <= 32'b01101110101010000001010001001001;
12'b010110100001: dataA <= 32'b00001110001101001011001010111001;
12'b010110100010: dataA <= 32'b00111000110010100001011101000110;
12'b010110100011: dataA <= 32'b00001011000010111000011110101011;
12'b010110100100: dataA <= 32'b10011101010011011001100000101110;
12'b010110100101: dataA <= 32'b00001101100110111000100110011100;
12'b010110100110: dataA <= 32'b11011010110101111101101000011110;
12'b010110100111: dataA <= 32'b00000100011010110101100010111010;
12'b010110101000: dataA <= 32'b11001110101010110001000100100110;
12'b010110101001: dataA <= 32'b00000101110110001101011111100001;
12'b010110101010: dataA <= 32'b10011010110001101110001001010111;
12'b010110101011: dataA <= 32'b00000010001110101000110100100001;
12'b010110101100: dataA <= 32'b01110100101001010100111000010010;
12'b010110101101: dataA <= 32'b00000111001110100110110100001011;
12'b010110101110: dataA <= 32'b11100000111111010001010111101010;
12'b010110101111: dataA <= 32'b00001001011000011101110101011011;
12'b010110110000: dataA <= 32'b00101101000011000011000100001110;
12'b010110110001: dataA <= 32'b00001000000100010100011110001100;
12'b010110110010: dataA <= 32'b10100011110001010011001010101100;
12'b010110110011: dataA <= 32'b00000010100100001110101101100110;
12'b010110110100: dataA <= 32'b01101100011001010000010110001001;
12'b010110110101: dataA <= 32'b00001000000001011110100110001001;
12'b010110110110: dataA <= 32'b01011000110001000010001000000111;
12'b010110110111: dataA <= 32'b00001000011000010101110111011001;
12'b010110111000: dataA <= 32'b00111011011110100100001101001111;
12'b010110111001: dataA <= 32'b00001101111010101101101111010110;
12'b010110111010: dataA <= 32'b10101011001000110001000011101011;
12'b010110111011: dataA <= 32'b00001011111101100011110110000100;
12'b010110111100: dataA <= 32'b01110000001111000100011111010001;
12'b010110111101: dataA <= 32'b00000110101011010000111010010000;
12'b010110111110: dataA <= 32'b10010001110011001011100011010101;
12'b010110111111: dataA <= 32'b00001010010011011111011101000110;
12'b010111000000: dataA <= 32'b10011110111101110010011010001001;
12'b010111000001: dataA <= 32'b00001100000011000100101010011010;
12'b010111000010: dataA <= 32'b00001000111111011100111011110110;
12'b010111000011: dataA <= 32'b00001110001011101110110100001011;
12'b010111000100: dataA <= 32'b11001111001000110010000000101101;
12'b010111000101: dataA <= 32'b00001011000010100100011101100011;
12'b010111000110: dataA <= 32'b10011001111001111000011010100011;
12'b010111000111: dataA <= 32'b00001011010110100111110011110100;
12'b010111001000: dataA <= 32'b10100110110001000011001100001010;
12'b010111001001: dataA <= 32'b00000111011101100111110011000010;
12'b010111001010: dataA <= 32'b00100111100000101001011011100111;
12'b010111001011: dataA <= 32'b00000000110100101011000010111101;
12'b010111001100: dataA <= 32'b00001101000010110011101001010010;
12'b010111001101: dataA <= 32'b00001110110001111011010111001010;
12'b010111001110: dataA <= 32'b10110111100101100110101100010110;
12'b010111001111: dataA <= 32'b00000111000001010110011110110101;
12'b010111010000: dataA <= 32'b01011001100001001000100111001001;
12'b010111010001: dataA <= 32'b00000111111110010101110110000101;
12'b010111010010: dataA <= 32'b01101010110000010010001001001110;
12'b010111010011: dataA <= 32'b00001110101110011101010001111011;
12'b010111010100: dataA <= 32'b01110000111000110001000110000111;
12'b010111010101: dataA <= 32'b00000111011011111011011101101100;
12'b010111010110: dataA <= 32'b10111010100100100011011101000111;
12'b010111010111: dataA <= 32'b00001010001010001110111101100011;
12'b010111011000: dataA <= 32'b11000011001110110100100011011011;
12'b010111011001: dataA <= 32'b00001000101000101100011110111010;
12'b010111011010: dataA <= 32'b00101111100101010010000011001011;
12'b010111011011: dataA <= 32'b00000011110111010001110010101101;
12'b010111011100: dataA <= 32'b01001101101111000001111010001010;
12'b010111011101: dataA <= 32'b00000011101100100000101101011110;
12'b010111011110: dataA <= 32'b00111011000111001101011111010100;
12'b010111011111: dataA <= 32'b00001100100100101010011010011101;
12'b010111100000: dataA <= 32'b01100100001110100011110111110010;
12'b010111100001: dataA <= 32'b00000110110110110111101010100000;
12'b010111100010: dataA <= 32'b10010011001011101100010010111011;
12'b010111100011: dataA <= 32'b00000100110001011101000100001100;
12'b010111100100: dataA <= 32'b10101111000110011100010100010111;
12'b010111100101: dataA <= 32'b00000110101000010010101111110011;
12'b010111100110: dataA <= 32'b10100101000110001001110110101100;
12'b010111100111: dataA <= 32'b00000001001000111010100111011010;
12'b010111101000: dataA <= 32'b01010010101001111100011110101111;
12'b010111101001: dataA <= 32'b00001010101001100000101110100000;
12'b010111101010: dataA <= 32'b00001111101010001101101010110101;
12'b010111101011: dataA <= 32'b00001101011010011101111011001101;
12'b010111101100: dataA <= 32'b00111010100110101001011000000111;
12'b010111101101: dataA <= 32'b00001000011010101011100100111100;
12'b010111101110: dataA <= 32'b10101110111000001101011110101110;
12'b010111101111: dataA <= 32'b00001100011100111001100000111100;
12'b010111110000: dataA <= 32'b11010111010110001100111111010100;
12'b010111110001: dataA <= 32'b00001011101111000111011111010011;
12'b010111110010: dataA <= 32'b01100100011100110001000001001000;
12'b010111110011: dataA <= 32'b00000100110010000011010101101000;
12'b010111110100: dataA <= 32'b11011011100111001100111001110110;
12'b010111110101: dataA <= 32'b00000110010101100101010011010100;
12'b010111110110: dataA <= 32'b11101100100001110001100000101100;
12'b010111110111: dataA <= 32'b00001110001011001011010010101000;
12'b010111111000: dataA <= 32'b11110110101010010001001100000101;
12'b010111111001: dataA <= 32'b00001001100001110100010110100010;
12'b010111111010: dataA <= 32'b01011111010011001001000000110001;
12'b010111111011: dataA <= 32'b00001100100100110100011110011100;
12'b010111111100: dataA <= 32'b01011010110110000101101001111110;
12'b010111111101: dataA <= 32'b00000101011100111001011010110010;
12'b010111111110: dataA <= 32'b01001100110010100000110011101000;
12'b010111111111: dataA <= 32'b00000110010111010001100111010001;
12'b011000000000: dataA <= 32'b00011000110001111110001010010111;
12'b011000000001: dataA <= 32'b00000010010000101000110000010010;
12'b011000000010: dataA <= 32'b00110010100001011101001000010010;
12'b011000000011: dataA <= 32'b00000111001110100110110000001100;
12'b011000000100: dataA <= 32'b00100000111111000000110111001010;
12'b011000000101: dataA <= 32'b00001010011000100001110101011100;
12'b011000000110: dataA <= 32'b00101100111110111010100100010000;
12'b011000000111: dataA <= 32'b00000111000100010000100010001100;
12'b011000001000: dataA <= 32'b11100111110001010011011010001011;
12'b011000001001: dataA <= 32'b00000010000110001100110101110110;
12'b011000001010: dataA <= 32'b01101000010101000000110101101010;
12'b011000001011: dataA <= 32'b00000110100001011010100101111001;
12'b011000001100: dataA <= 32'b11011000110100111010100111000111;
12'b011000001101: dataA <= 32'b00001001010111011011110111000000;
12'b011000001110: dataA <= 32'b01111101010010100011111100101101;
12'b011000001111: dataA <= 32'b00001110010111110001101011100101;
12'b011000010000: dataA <= 32'b10101101000100100001100011001101;
12'b011000010001: dataA <= 32'b00001100111011101001110010001100;
12'b011000010010: dataA <= 32'b01101010001011000011111111001111;
12'b011000010011: dataA <= 32'b00000110001100001110111101111000;
12'b011000010100: dataA <= 32'b11010101111011001011000011110110;
12'b011000010101: dataA <= 32'b00001010110010100001011101010110;
12'b011000010110: dataA <= 32'b10011110111101101010011001001000;
12'b011000010111: dataA <= 32'b00001010100010000100110110010010;
12'b011000011000: dataA <= 32'b11001001000111100100011100010100;
12'b011000011001: dataA <= 32'b00001101001000101110110000001011;
12'b011000011010: dataA <= 32'b00010001010000101010100000110000;
12'b011000011011: dataA <= 32'b00001001100001100010011101100100;
12'b011000011100: dataA <= 32'b11011111111001100000011001100010;
12'b011000011101: dataA <= 32'b00001011110101101101101111110011;
12'b011000011110: dataA <= 32'b00100100110001000011101011101000;
12'b011000011111: dataA <= 32'b00001000111101101101101110111010;
12'b011000100000: dataA <= 32'b11101011011100011001111010100101;
12'b011000100001: dataA <= 32'b00000001010111101010111111000100;
12'b011000100010: dataA <= 32'b10001111001010110011011001110001;
12'b011000100011: dataA <= 32'b00001110101110111101001110111001;
12'b011000100100: dataA <= 32'b01111011011101110110101100110101;
12'b011000100101: dataA <= 32'b00000101100001010010100010111101;
12'b011000100110: dataA <= 32'b00011101100100111000110110101001;
12'b011000100111: dataA <= 32'b00001001011110011001111010001101;
12'b011000101000: dataA <= 32'b01101000101100001010111001001101;
12'b011000101001: dataA <= 32'b00001110001011011111010001110011;
12'b011000101010: dataA <= 32'b10110000110000100001100101001000;
12'b011000101011: dataA <= 32'b00001000011011111101010001101100;
12'b011000101100: dataA <= 32'b11111000011100100011111100100101;
12'b011000101101: dataA <= 32'b00001001101001001111000101100011;
12'b011000101110: dataA <= 32'b10000101011010111100000100111101;
12'b011000101111: dataA <= 32'b00001000000111101010011010110010;
12'b011000110000: dataA <= 32'b11110011011101001010010010101101;
12'b011000110001: dataA <= 32'b00000100111001010111111010110100;
12'b011000110010: dataA <= 32'b10010001110110110001011001101001;
12'b011000110011: dataA <= 32'b00000011001110011110101101101110;
12'b011000110100: dataA <= 32'b11111010111011010100111111010001;
12'b011000110101: dataA <= 32'b00001011000010100110010110100100;
12'b011000110110: dataA <= 32'b01100000001110011011101000010010;
12'b011000110111: dataA <= 32'b00000111110111111001011110010000;
12'b011000111000: dataA <= 32'b01010011001111101011100100011100;
12'b011000111001: dataA <= 32'b00000100110010011101000100001101;
12'b011000111010: dataA <= 32'b11110001000010100100010101011000;
12'b011000111011: dataA <= 32'b00000110001000010000110111110010;
12'b011000111100: dataA <= 32'b00100101000001111001110110101100;
12'b011000111101: dataA <= 32'b00000000101011111000011111010010;
12'b011000111110: dataA <= 32'b01010000110001111100011110001100;
12'b011000111111: dataA <= 32'b00001001101000011110101110010000;
12'b011001000000: dataA <= 32'b10010101110010010101101011010100;
12'b011001000001: dataA <= 32'b00001110011000100001111011010100;
12'b011001000010: dataA <= 32'b10111000011110010001000111000111;
12'b011001000011: dataA <= 32'b00001001011010101101100001000100;
12'b011001000100: dataA <= 32'b00101110110100011101111110001011;
12'b011001000101: dataA <= 32'b00001101011010111011010101000101;
12'b011001000110: dataA <= 32'b01011001011010001100111111010001;
12'b011001000111: dataA <= 32'b00001011101110001011101011010011;
12'b011001001000: dataA <= 32'b01100010011100100001100000101011;
12'b011001001001: dataA <= 32'b00000100110011000111011101010000;
12'b011001001010: dataA <= 32'b01011111100111001100011010110101;
12'b011001001011: dataA <= 32'b00000110110101100111001111010100;
12'b011001001100: dataA <= 32'b10101000011101100001100000101111;
12'b011001001101: dataA <= 32'b00001101001000001101011010011000;
12'b011001001110: dataA <= 32'b10110100100010000001001010100011;
12'b011001001111: dataA <= 32'b00001000000001110000001110011010;
12'b011001010000: dataA <= 32'b01100001010010111000110000110100;
12'b011001010001: dataA <= 32'b00001011100010110010010110100100;
12'b011001010010: dataA <= 32'b00011000111010001101011011011101;
12'b011001010011: dataA <= 32'b00000110011101111011010010101010;
12'b011001010100: dataA <= 32'b11001100111010001000100010101010;
12'b011001010101: dataA <= 32'b00000111010111010101101011000000;
12'b011001010110: dataA <= 32'b11011000110110001110001010110110;
12'b011001010111: dataA <= 32'b00000010010010100110101100001010;
12'b011001011000: dataA <= 32'b11101110011101100101011000110010;
12'b011001011001: dataA <= 32'b00000111001110100100110000001100;
12'b011001011010: dataA <= 32'b01100000111110101000100110101010;
12'b011001011011: dataA <= 32'b00001011010110100111110001100100;
12'b011001011100: dataA <= 32'b00101010111010110010010100010001;
12'b011001011101: dataA <= 32'b00000110000101001110101010001100;
12'b011001011110: dataA <= 32'b11101101101101001011101001101010;
12'b011001011111: dataA <= 32'b00000001001001001100111110000110;
12'b011001100000: dataA <= 32'b10100010010000101001010101001011;
12'b011001100001: dataA <= 32'b00000101000001011000100101101001;
12'b011001100010: dataA <= 32'b10010110111000110011000110100111;
12'b011001100011: dataA <= 32'b00001001110111100001111010110000;
12'b011001100100: dataA <= 32'b11111101000110100011111100001011;
12'b011001100101: dataA <= 32'b00001111010101110101100011101100;
12'b011001100110: dataA <= 32'b10101100111100010010000011001111;
12'b011001100111: dataA <= 32'b00001101111001101101101110001100;
12'b011001101000: dataA <= 32'b01100100000111000011101110101100;
12'b011001101001: dataA <= 32'b00000110001100010001000101101000;
12'b011001101010: dataA <= 32'b00011011111011000010100100011000;
12'b011001101011: dataA <= 32'b00001010110001100101011101101111;
12'b011001101100: dataA <= 32'b01011110111101100010011000101000;
12'b011001101101: dataA <= 32'b00001001000001000011000010001010;
12'b011001101110: dataA <= 32'b10001001001111100011111100010011;
12'b011001101111: dataA <= 32'b00001100100110101100101000001100;
12'b011001110000: dataA <= 32'b01010011010100100011000000110010;
12'b011001110001: dataA <= 32'b00001000000001011110011101101100;
12'b011001110010: dataA <= 32'b01100101111001001000101000000010;
12'b011001110011: dataA <= 32'b00001100010011110001101011110011;
12'b011001110100: dataA <= 32'b11100010101101000011111010100111;
12'b011001110101: dataA <= 32'b00001010011101110001101010101001;
12'b011001110110: dataA <= 32'b01101101011000010010101001100101;
12'b011001110111: dataA <= 32'b00000010011001101010111011001100;
12'b011001111000: dataA <= 32'b01001111010010110011001001110001;
12'b011001111001: dataA <= 32'b00001110101011111101000010101001;
12'b011001111010: dataA <= 32'b11111101010010001110101101010011;
12'b011001111011: dataA <= 32'b00000100000010010000100111000100;
12'b011001111100: dataA <= 32'b00011111100100101001010110001001;
12'b011001111101: dataA <= 32'b00001010111110011111111010010101;
12'b011001111110: dataA <= 32'b01100110101000001011101000101101;
12'b011001111111: dataA <= 32'b00001101101001100001010001110011;
12'b011010000000: dataA <= 32'b10101110101100010010000100101001;
12'b011010000001: dataA <= 32'b00001001011010111101000101110100;
12'b011010000010: dataA <= 32'b00110100010100100100011011000011;
12'b011010000011: dataA <= 32'b00001001001001001111001001100100;
12'b011010000100: dataA <= 32'b01000111100010111011110110011110;
12'b011010000101: dataA <= 32'b00000111001000100110010110100010;
12'b011010000110: dataA <= 32'b10110101010100111010100010101111;
12'b011010000111: dataA <= 32'b00000101111010011011111010110100;
12'b011010001000: dataA <= 32'b10010111111010100001001001001001;
12'b011010001001: dataA <= 32'b00000011001111011110101101111110;
12'b011010001010: dataA <= 32'b10111010101111011100011111001110;
12'b011010001011: dataA <= 32'b00001010000001100010010010100100;
12'b011010001100: dataA <= 32'b01011010001110011011101000010010;
12'b011010001101: dataA <= 32'b00001000010111111101010101111000;
12'b011010001110: dataA <= 32'b11010101010011101010110101011110;
12'b011010001111: dataA <= 32'b00000100110011011111001000011101;
12'b011010010000: dataA <= 32'b00101110111010100100000110011001;
12'b011010010001: dataA <= 32'b00000101001001010000111011101010;
12'b011010010010: dataA <= 32'b10100101000001110001110110001101;
12'b011010010011: dataA <= 32'b00000000101110110100010111000001;
12'b011010010100: dataA <= 32'b01001110110101111100011101101010;
12'b011010010101: dataA <= 32'b00001001000111011110101101111000;
12'b011010010110: dataA <= 32'b00011001110110011101101011110010;
12'b011010010111: dataA <= 32'b00001110110101100111110111010100;
12'b011010011000: dataA <= 32'b11110100010110000000110110100111;
12'b011010011001: dataA <= 32'b00001010011001110001011101000100;
12'b011010011010: dataA <= 32'b01101100101100101110101101101001;
12'b011010011011: dataA <= 32'b00001110010111111101001001001101;
12'b011010011100: dataA <= 32'b11011011011010010100111111001110;
12'b011010011101: dataA <= 32'b00001011001101001111110011001010;
12'b011010011110: dataA <= 32'b11011110011100010010000000101110;
12'b011010011111: dataA <= 32'b00000101010100001011101001000000;
12'b011010100000: dataA <= 32'b10100011100111001011111010110100;
12'b011010100001: dataA <= 32'b00000111010110100111001111010011;
12'b011010100010: dataA <= 32'b10100110011101010001110000110010;
12'b011010100011: dataA <= 32'b00001100100110010001011110000000;
12'b011010100100: dataA <= 32'b01110000011001110001001001100010;
12'b011010100101: dataA <= 32'b00000110100001101010001010010010;
12'b011010100110: dataA <= 32'b00100001010010100000010001010111;
12'b011010100111: dataA <= 32'b00001010000001101100001110100100;
12'b011010101000: dataA <= 32'b11011000111010011101011100011100;
12'b011010101001: dataA <= 32'b00000111111101111101000110011001;
12'b011010101010: dataA <= 32'b10001101000001111000100010101100;
12'b011010101011: dataA <= 32'b00000111110111011001101110101000;
12'b011010101100: dataA <= 32'b10010110111010010110001011010100;
12'b011010101101: dataA <= 32'b00000010110100100100101100001011;
12'b011010101110: dataA <= 32'b10101010010101101101101000110010;
12'b011010101111: dataA <= 32'b00000110101111100010101100010101;
12'b011010110000: dataA <= 32'b01100000111110010000010110001011;
12'b011010110001: dataA <= 32'b00001011110101101011101101100100;
12'b011010110010: dataA <= 32'b00101010110010101001110100110010;
12'b011010110011: dataA <= 32'b00000101000110001100110010001100;
12'b011010110100: dataA <= 32'b10110001101001001100001001001001;
12'b011010110101: dataA <= 32'b00000000101100001101000110010110;
12'b011010110110: dataA <= 32'b11011110010000011001110100101100;
12'b011010110111: dataA <= 32'b00000100000011010110101001011001;
12'b011010111000: dataA <= 32'b01010110111100101011100101101000;
12'b011010111001: dataA <= 32'b00001010010110100101110110011000;
12'b011010111010: dataA <= 32'b00111100111010100011101011101001;
12'b011010111011: dataA <= 32'b00001111010010110111010111101100;
12'b011010111100: dataA <= 32'b01101100111000001010110011010000;
12'b011010111101: dataA <= 32'b00001110110111110001100110010100;
12'b011010111110: dataA <= 32'b10011110000111000011001110001001;
12'b011010111111: dataA <= 32'b00000101101101010001001001010000;
12'b011011000000: dataA <= 32'b00100001111010111010000101011001;
12'b011011000001: dataA <= 32'b00001010110000100111011001111111;
12'b011011000010: dataA <= 32'b01011110111101011010100111101000;
12'b011011000011: dataA <= 32'b00000111100001000101001010000010;
12'b011011000100: dataA <= 32'b01001011010111011011001100110001;
12'b011011000101: dataA <= 32'b00001011100101101010100100001101;
12'b011011000110: dataA <= 32'b01010101011000011011110001010101;
12'b011011000111: dataA <= 32'b00000110100001011010011101101100;
12'b011011001000: dataA <= 32'b10101001111000111000110110100010;
12'b011011001001: dataA <= 32'b00001100010001110101100011101010;
12'b011011001010: dataA <= 32'b10100000101101000100011010000110;
12'b011011001011: dataA <= 32'b00001011011100110101100010100001;
12'b011011001100: dataA <= 32'b11101111010000001011011000100100;
12'b011011001101: dataA <= 32'b00000011011011101000110111001011;
12'b011011001110: dataA <= 32'b00010001010110101010111001110000;
12'b011011001111: dataA <= 32'b00001110001001111100110110011001;
12'b011011010000: dataA <= 32'b01111101000110011110101101010001;
12'b011011010001: dataA <= 32'b00000011000100001110101111000100;
12'b011011010010: dataA <= 32'b11100011100100011010000101101010;
12'b011011010011: dataA <= 32'b00001011111100100101111010011100;
12'b011011010100: dataA <= 32'b10100100101000001100011000101101;
12'b011011010101: dataA <= 32'b00001100100111100011010001101011;
12'b011011010110: dataA <= 32'b10101100100100001010110100001011;
12'b011011010111: dataA <= 32'b00001010011010111100111001110100;
12'b011011011000: dataA <= 32'b01101110001100101100111010000010;
12'b011011011001: dataA <= 32'b00001000001000010001010001100100;
12'b011011011010: dataA <= 32'b00001011101010110011010111111110;
12'b011011011011: dataA <= 32'b00000110101000100010010110011010;
12'b011011011100: dataA <= 32'b00110111001100111011000010110001;
12'b011011011101: dataA <= 32'b00000110111010100001111010111100;
12'b011011011110: dataA <= 32'b10011101111010010000111000001000;
12'b011011011111: dataA <= 32'b00000011010001011100101110001110;
12'b011011100000: dataA <= 32'b01111000100111011011101111001011;
12'b011011100001: dataA <= 32'b00001000100001011100010010101100;
12'b011011100010: dataA <= 32'b01010110010010011011011000010010;
12'b011011100011: dataA <= 32'b00001001010110111101001001100000;
12'b011011100100: dataA <= 32'b10010111010111100010010110111110;
12'b011011100101: dataA <= 32'b00000101010100011111001000101110;
12'b011011100110: dataA <= 32'b10101110110110100011110111011010;
12'b011011100111: dataA <= 32'b00000100101010010001000011011001;
12'b011011101000: dataA <= 32'b00100100111101100001110110001110;
12'b011011101001: dataA <= 32'b00000000110001101110001110110001;
12'b011011101010: dataA <= 32'b01001110111110000100011101000111;
12'b011011101011: dataA <= 32'b00001000000111011100101101100000;
12'b011011101100: dataA <= 32'b10011111110110100101011011110001;
12'b011011101101: dataA <= 32'b00001111010010101101110011010011;
12'b011011101110: dataA <= 32'b00101110001101110001000101101000;
12'b011011101111: dataA <= 32'b00001010111000110011010101001101;
12'b011011110000: dataA <= 32'b10101010101000111111001100100111;
12'b011011110001: dataA <= 32'b00001111010101111100111101010101;
12'b011011110010: dataA <= 32'b10011111011110011100101111001011;
12'b011011110011: dataA <= 32'b00001010101011010011110111000010;
12'b011011110100: dataA <= 32'b01011010011100001010110000110001;
12'b011011110101: dataA <= 32'b00000101110101001111110000101001;
12'b011011110110: dataA <= 32'b00100111100011001011011011010010;
12'b011011110111: dataA <= 32'b00000111110110101001001011010011;
12'b011011111000: dataA <= 32'b10100010011001000010000000110101;
12'b011011111001: dataA <= 32'b00001011100101010011100101101000;
12'b011011111010: dataA <= 32'b01101100010001100001011000000010;
12'b011011111011: dataA <= 32'b00000101000001100100000110001010;
12'b011011111100: dataA <= 32'b11100011010010010000010010011001;
12'b011011111101: dataA <= 32'b00001000100001101000001010100011;
12'b011011111110: dataA <= 32'b11011000111110100101001101011010;
12'b011011111111: dataA <= 32'b00001001011101111100111010001001;
12'b011100000000: dataA <= 32'b01001101001001100000100010001110;
12'b011100000001: dataA <= 32'b00001000110111011111110010010000;
12'b011100000010: dataA <= 32'b01010110111110100101111011110011;
12'b011100000011: dataA <= 32'b00000011010110100010101000001100;
12'b011100000100: dataA <= 32'b00100110010001110101101001010001;
12'b011100000101: dataA <= 32'b00000110101111100000101100011110;
12'b011100000110: dataA <= 32'b10100000111101111000010101101100;
12'b011100000111: dataA <= 32'b00001100010100110001101001100100;
12'b011100001000: dataA <= 32'b11101000101110011001110101010100;
12'b011100001001: dataA <= 32'b00000100000111001010111010001011;
12'b011100001010: dataA <= 32'b10110101100001001100011000101001;
12'b011100001011: dataA <= 32'b00000000101111001111001110100110;
12'b011100001100: dataA <= 32'b00011010010000010010010100001101;
12'b011100001101: dataA <= 32'b00000010100101010100101101001010;
12'b011100001110: dataA <= 32'b01010110111100101100000101001001;
12'b011100001111: dataA <= 32'b00001011010101101011110110000000;
12'b011100010000: dataA <= 32'b10111100101110011011011011001000;
12'b011100010001: dataA <= 32'b00001111001111111001001111101011;
12'b011100010010: dataA <= 32'b01101010110100001011100011010010;
12'b011100010011: dataA <= 32'b00001111010100110101011110010100;
12'b011100010100: dataA <= 32'b11011000000110111010101101100111;
12'b011100010101: dataA <= 32'b00000101101110010011010000111000;
12'b011100010110: dataA <= 32'b00100111111010101001110110011010;
12'b011100010111: dataA <= 32'b00001010101111101001010110010111;
12'b011100011000: dataA <= 32'b01011110111101010010110111001000;
12'b011100011001: dataA <= 32'b00000110000001000101010101110010;
12'b011100011010: dataA <= 32'b11001111011111010010101100101111;
12'b011100011011: dataA <= 32'b00001010100100100110100000011101;
12'b011100011100: dataA <= 32'b10010111011100011100010001111000;
12'b011100011101: dataA <= 32'b00000101100001011000100001101100;
12'b011100011110: dataA <= 32'b11101111110000101001010101100011;
12'b011100011111: dataA <= 32'b00001100010000110111011011100001;
12'b011100100000: dataA <= 32'b01100000101101000100101001000101;
12'b011100100001: dataA <= 32'b00001100111010110111011010010001;
12'b011100100010: dataA <= 32'b10110001001100001011110111100100;
12'b011100100011: dataA <= 32'b00000100011101101000110011001011;
12'b011100100100: dataA <= 32'b11010011011010100010101001101111;
12'b011100100101: dataA <= 32'b00001101000110111010101010000000;
12'b011100100110: dataA <= 32'b00111100111010101110011101001110;
12'b011100100111: dataA <= 32'b00000010000110001100110111000100;
12'b011100101000: dataA <= 32'b11100111100000001010100101001011;
12'b011100101001: dataA <= 32'b00001101011010101011110110011100;
12'b011100101010: dataA <= 32'b10100010100100001101001000001100;
12'b011100101011: dataA <= 32'b00001011100101100101010001101011;
12'b011100101100: dataA <= 32'b11101010100000001011100011101100;
12'b011100101101: dataA <= 32'b00001011011001111100101101111100;
12'b011100101110: dataA <= 32'b01101010000100101101011000100010;
12'b011100101111: dataA <= 32'b00000111101000010011010101100100;
12'b011100110000: dataA <= 32'b00010001110010110011001001011110;
12'b011100110001: dataA <= 32'b00000101101001011100010110010010;
12'b011100110010: dataA <= 32'b11111001000000110011100011010011;
12'b011100110011: dataA <= 32'b00000111111011100111111010111011;
12'b011100110100: dataA <= 32'b01100011111001111000110111101000;
12'b011100110101: dataA <= 32'b00000011110011011010110010011110;
12'b011100110110: dataA <= 32'b00110100011011010011001110101001;
12'b011100110111: dataA <= 32'b00000111000001011000010110101100;
12'b011100111000: dataA <= 32'b10010010010110010011001000110001;
12'b011100111001: dataA <= 32'b00001001110110111100111101001000;
12'b011100111010: dataA <= 32'b00011001011011010001101000011110;
12'b011100111011: dataA <= 32'b00000101110101011111001000111111;
12'b011100111100: dataA <= 32'b00101100101110100011101000011010;
12'b011100111101: dataA <= 32'b00000100001100010001000111001001;
12'b011100111110: dataA <= 32'b11100100111101010010000110001110;
12'b011100111111: dataA <= 32'b00000000110100101010000110100000;
12'b011101000000: dataA <= 32'b10001111000110000100011100000101;
12'b011101000001: dataA <= 32'b00000111000111011010110001001000;
12'b011101000010: dataA <= 32'b00100011110110101101001100001111;
12'b011101000011: dataA <= 32'b00001111010000110001101111001011;
12'b011101000100: dataA <= 32'b10101010000101011001000101001001;
12'b011101000101: dataA <= 32'b00001011110111110101001101010101;
12'b011101000110: dataA <= 32'b11101000100101001111011011100101;
12'b011101000111: dataA <= 32'b00001111010010111100110001011101;
12'b011101001000: dataA <= 32'b00100001011110011100011110101001;
12'b011101001001: dataA <= 32'b00001010101010011001111010111010;
12'b011101001010: dataA <= 32'b11011000100000001011100000110100;
12'b011101001011: dataA <= 32'b00000110010110010011110100011001;
12'b011101001100: dataA <= 32'b10101001100011001010111011110001;
12'b011101001101: dataA <= 32'b00001000110110101001000111001010;
12'b011101001110: dataA <= 32'b11011110011000111010100001110111;
12'b011101001111: dataA <= 32'b00001010100100010111101001011000;
12'b011101010000: dataA <= 32'b01101000001101010001010111000010;
12'b011101010001: dataA <= 32'b00000100000011011110000110000010;
12'b011101010010: dataA <= 32'b10100101001101111000010011011011;
12'b011101010011: dataA <= 32'b00000111000001100010001010100011;
12'b011101010100: dataA <= 32'b11011001000010100100111110010111;
12'b011101010101: dataA <= 32'b00001010011100111010101110000001;
12'b011101010110: dataA <= 32'b01001101010001010000110010010000;
12'b011101010111: dataA <= 32'b00001001010111100011110010000000;
12'b011101011000: dataA <= 32'b00010110111110101101101011110010;
12'b011101011001: dataA <= 32'b00000100011000100000101000001101;
12'b011101011010: dataA <= 32'b10100010010001111101101001010001;
12'b011101011011: dataA <= 32'b00000110101111100000101100101110;
12'b011101011100: dataA <= 32'b11100000111101100000010101001101;
12'b011101011101: dataA <= 32'b00001100010010110101100001101100;
12'b011101011110: dataA <= 32'b11100110101110001001100101010101;
12'b011101011111: dataA <= 32'b00000011101001001011000010001011;
12'b011101100000: dataA <= 32'b01110111011001010100101000001001;
12'b011101100001: dataA <= 32'b00000000110010001111010010110110;
12'b011101100010: dataA <= 32'b01010110010100001011000100001111;
12'b011101100011: dataA <= 32'b00000001100111010010110001000010;
12'b011101100100: dataA <= 32'b01010111000000101100100100101010;
12'b011101100101: dataA <= 32'b00001011110100101111101101101000;
12'b011101100110: dataA <= 32'b11111010100010011011001010000111;
12'b011101100111: dataA <= 32'b00001111001100111011000011100010;
12'b011101101000: dataA <= 32'b00101010110000001100010011110100;
12'b011101101001: dataA <= 32'b00001111010001110111010110010100;
12'b011101101010: dataA <= 32'b01010100001010110010011100100101;
12'b011101101011: dataA <= 32'b00000101001111010101010100101001;
12'b011101101100: dataA <= 32'b11101101110110011001100111011011;
12'b011101101101: dataA <= 32'b00001010101110101011010010100110;
12'b011101101110: dataA <= 32'b10011110111101001011010110001000;
12'b011101101111: dataA <= 32'b00000101000010001001011101101010;
12'b011101110000: dataA <= 32'b10010001100111001010001100101101;
12'b011101110001: dataA <= 32'b00001001000011100100100000100110;
12'b011101110010: dataA <= 32'b10011011100000100100110010111010;
12'b011101110011: dataA <= 32'b00000100000011010100100101110100;
12'b011101110100: dataA <= 32'b01110011101100011010000100100100;
12'b011101110101: dataA <= 32'b00001100001110111001001111010001;
12'b011101110110: dataA <= 32'b01011110101101001101001000000101;
12'b011101110111: dataA <= 32'b00001101011000111001001110000001;
12'b011101111000: dataA <= 32'b00110001000100001100100110100100;
12'b011101111001: dataA <= 32'b00000101111110100110101111000011;
12'b011101111010: dataA <= 32'b00010111100010010010011001101110;
12'b011101111011: dataA <= 32'b00001100000101111000011101110001;
12'b011101111100: dataA <= 32'b10111100101110110110001101001100;
12'b011101111101: dataA <= 32'b00000001001000001010111111000011;
12'b011101111110: dataA <= 32'b10101001011100001011010100101101;
12'b011101111111: dataA <= 32'b00001110011000110001110010100100;
12'b011110000000: dataA <= 32'b11011110100100010101110111101100;
12'b011110000001: dataA <= 32'b00001010100100100101010001101011;
12'b011110000010: dataA <= 32'b11100110011100001100010011101110;
12'b011110000011: dataA <= 32'b00001100010111111010100010000100;
12'b011110000100: dataA <= 32'b10100100000100111101110111000010;
12'b011110000101: dataA <= 32'b00000110101001010101011001101100;
12'b011110000110: dataA <= 32'b11010101111010101010111010011110;
12'b011110000111: dataA <= 32'b00000101001010011000010110000001;
12'b011110001000: dataA <= 32'b01110110111000110100000011010101;
12'b011110001001: dataA <= 32'b00001000111011101101110110110011;
12'b011110001010: dataA <= 32'b01101001111001101000110110101001;
12'b011110001011: dataA <= 32'b00000100010100011000110010101110;
12'b011110001100: dataA <= 32'b11110000010111001010101101100110;
12'b011110001101: dataA <= 32'b00000101100001010100011010101011;
12'b011110001110: dataA <= 32'b00001110011110010011001000110001;
12'b011110001111: dataA <= 32'b00001010010101111100110000110001;
12'b011110010000: dataA <= 32'b01011011011011000001011001111110;
12'b011110010001: dataA <= 32'b00000110110110100001001001001111;
12'b011110010010: dataA <= 32'b10101010101010011011101001011010;
12'b011110010011: dataA <= 32'b00000100001101010001001110111000;
12'b011110010100: dataA <= 32'b10100100111001001010010101101111;
12'b011110010101: dataA <= 32'b00000001010111100100000110001000;
12'b011110010110: dataA <= 32'b00001111001010000100011011000100;
12'b011110010111: dataA <= 32'b00000110100111011000110000110001;
12'b011110011000: dataA <= 32'b10101001110010110100101011101110;
12'b011110011001: dataA <= 32'b00001111001101110101100111001010;
12'b011110011010: dataA <= 32'b11100100000101001001010100101010;
12'b011110011011: dataA <= 32'b00001100010101110111000101011101;
12'b011110011100: dataA <= 32'b00100110100001100111101010100100;
12'b011110011101: dataA <= 32'b00001111001111111010101001101110;
12'b011110011110: dataA <= 32'b11100101011010011100011101100110;
12'b011110011111: dataA <= 32'b00001001101001011111111010101001;
12'b011110100000: dataA <= 32'b01010100100100001100010001010111;
12'b011110100001: dataA <= 32'b00000110110110011001111000010010;
12'b011110100010: dataA <= 32'b01101101011111000010101011110000;
12'b011110100011: dataA <= 32'b00001001010101101011000011000010;
12'b011110100100: dataA <= 32'b00011010011000110011000010011010;
12'b011110100101: dataA <= 32'b00001001000011011011101001001001;
12'b011110100110: dataA <= 32'b01100010001001000001110101100011;
12'b011110100111: dataA <= 32'b00000010100100011010000101110010;
12'b011110101000: dataA <= 32'b10100111001101100000010100011101;
12'b011110101001: dataA <= 32'b00000101100001011100001010011011;
12'b011110101010: dataA <= 32'b11011001000110101100101111010101;
12'b011110101011: dataA <= 32'b00001011011011111000100101110001;
12'b011110101100: dataA <= 32'b01001111010100111001010010010010;
12'b011110101101: dataA <= 32'b00001010010110100111101101101000;
12'b011110101110: dataA <= 32'b11010111000010110101011100010000;
12'b011110101111: dataA <= 32'b00000100111001011110101000010101;
12'b011110110000: dataA <= 32'b00011110010010001101101001010000;
12'b011110110001: dataA <= 32'b00000110110000011110101101000111;
12'b011110110010: dataA <= 32'b11100000111101010000100101001110;
12'b011110110011: dataA <= 32'b00001100110000110111011001101100;
12'b011110110100: dataA <= 32'b11100100101001111001100110010110;
12'b011110110101: dataA <= 32'b00000011001010001011001010001011;
12'b011110110110: dataA <= 32'b11111001001101010100110111001001;
12'b011110110111: dataA <= 32'b00000000110100010001011011000101;
12'b011110111000: dataA <= 32'b11010010011000001011110100010000;
12'b011110111001: dataA <= 32'b00000001001001010010110100111010;
12'b011110111010: dataA <= 32'b01010111000100110101000100001100;
12'b011110111011: dataA <= 32'b00001011110010110101101001011000;
12'b011110111100: dataA <= 32'b01110110011010010011001001000110;
12'b011110111101: dataA <= 32'b00001110101001111010111011011010;
12'b011110111110: dataA <= 32'b00101000101100001101000100010110;
12'b011110111111: dataA <= 32'b00001111001110111001001110010100;
12'b011111000000: dataA <= 32'b11001110001110100010001011100011;
12'b011111000001: dataA <= 32'b00000101010000010111011000011001;
12'b011111000010: dataA <= 32'b10110001110010001001101000011011;
12'b011111000011: dataA <= 32'b00001010101101101101001110110110;
12'b011111000100: dataA <= 32'b10011110111101001011100101101001;
12'b011111000101: dataA <= 32'b00000011100011001011101001100010;
12'b011111000110: dataA <= 32'b00010101101010111001101100001011;
12'b011111000111: dataA <= 32'b00001000000010100000100000111111;
12'b011111001000: dataA <= 32'b10011111100000101101010011111100;
12'b011111001001: dataA <= 32'b00000011000100010010101001110100;
12'b011111001010: dataA <= 32'b11110111100100001010100011000110;
12'b011111001011: dataA <= 32'b00001100001100111001000111000000;
12'b011111001100: dataA <= 32'b01011100101101010101010110100101;
12'b011111001101: dataA <= 32'b00001110010110111001000101101001;
12'b011111001110: dataA <= 32'b10110010111100010101010101100101;
12'b011111001111: dataA <= 32'b00000111011110100100101110111010;
12'b011111010000: dataA <= 32'b00011011100010001010011001101110;
12'b011111010001: dataA <= 32'b00001011000011110100010101100001;
12'b011111010010: dataA <= 32'b00111010100011000101101100101010;
12'b011111010011: dataA <= 32'b00000000101011001011000111000011;
12'b011111010100: dataA <= 32'b01101101011000001100000100101110;
12'b011111010101: dataA <= 32'b00001110110110110101101010100100;
12'b011111010110: dataA <= 32'b11011100100100100110010111101100;
12'b011111010111: dataA <= 32'b00001001100011100111001101101011;
12'b011111011000: dataA <= 32'b11100010011100001101000011010000;
12'b011111011001: dataA <= 32'b00001100110101110110011010000100;
12'b011111011010: dataA <= 32'b10011110000101001110010110000010;
12'b011111011011: dataA <= 32'b00000110001001011001011101101100;
12'b011111011100: dataA <= 32'b11011011111010100010101011111100;
12'b011111011101: dataA <= 32'b00000100101011010100011001110001;
12'b011111011110: dataA <= 32'b00110110110000110100100100010111;
12'b011111011111: dataA <= 32'b00001001111010110001101110110011;
12'b011111100000: dataA <= 32'b11101111110101011001000110001001;
12'b011111100001: dataA <= 32'b00000100110110011000110110111101;
12'b011111100010: dataA <= 32'b10101100001111000010001100100100;
12'b011111100011: dataA <= 32'b00000100000010010000011110101011;
12'b011111100100: dataA <= 32'b01001010100010001011001000110001;
12'b011111100101: dataA <= 32'b00001010110100111010100100100001;
12'b011111100110: dataA <= 32'b10011111011010110000111011011101;
12'b011111100111: dataA <= 32'b00000111010110100001001001100111;
12'b011111101000: dataA <= 32'b01101000100110011011011010011001;
12'b011111101001: dataA <= 32'b00000100001111010011010010100000;
12'b011111101010: dataA <= 32'b10100100111001000010110101110000;
12'b011111101011: dataA <= 32'b00000010011001011110000101111000;
12'b011111101100: dataA <= 32'b01010001010010000100011010000011;
12'b011111101101: dataA <= 32'b00000101101000011000110100100001;
12'b011111101110: dataA <= 32'b00101101101110110100011011101100;
12'b011111101111: dataA <= 32'b00001110101010111001011110111010;
12'b011111110000: dataA <= 32'b11011110000100111001110100001100;
12'b011111110001: dataA <= 32'b00001100110011110110111101101101;
12'b011111110010: dataA <= 32'b00100010100001111111101001100011;
12'b011111110011: dataA <= 32'b00001111001100111000011101111110;
12'b011111110100: dataA <= 32'b10100111011010011100001100100100;
12'b011111110101: dataA <= 32'b00001001001001100101111010011001;
12'b011111110110: dataA <= 32'b00010010101000001101000010011001;
12'b011111110111: dataA <= 32'b00000111110110011111111000001011;
12'b011111111000: dataA <= 32'b11101111010110110010001011101110;
12'b011111111001: dataA <= 32'b00001001110101101010111110110001;
12'b011111111010: dataA <= 32'b10010110011100110011100011111100;
12'b011111111011: dataA <= 32'b00001000000010011111101100110001;
12'b011111111100: dataA <= 32'b01011110001000110010010100100100;
12'b011111111101: dataA <= 32'b00000001100111010100001001101010;
12'b011111111110: dataA <= 32'b01100111001001001000100101111110;
12'b011111111111: dataA <= 32'b00000100000010011000001010011011;
12'b100000000000: dataA <= 32'b11011001000110101100011111010010;
12'b100000000001: dataA <= 32'b00001100111001110100011101100001;
12'b100000000010: dataA <= 32'b10010011011100101001100010110100;
12'b100000000011: dataA <= 32'b00001010110101101011101001010000;
12'b100000000100: dataA <= 32'b01010111000110111100111100001110;
12'b100000000101: dataA <= 32'b00000101111010011100101000100110;
12'b100000000110: dataA <= 32'b10011010010010010101101001010000;
12'b100000000111: dataA <= 32'b00000110110000011100101101010111;
12'b100000001000: dataA <= 32'b11100000111100111000110101001111;
12'b100000001001: dataA <= 32'b00001100101110111001010001110100;
12'b100000001010: dataA <= 32'b11100010101001101001100110110110;
12'b100000001011: dataA <= 32'b00000010101100001101010010001011;
12'b100000001100: dataA <= 32'b01111001000101011101000110101001;
12'b100000001101: dataA <= 32'b00000001110111010101011111001101;
12'b100000001110: dataA <= 32'b01001110100000001100100100010010;
12'b100000001111: dataA <= 32'b00000000101100010010111100110011;
12'b100000010000: dataA <= 32'b00100011010010100110010110010111;
12'b100000010001: dataA <= 32'b00001001001000110100010100001101;
12'b100000010010: dataA <= 32'b00001100010001100011010011001101;
12'b100000010011: dataA <= 32'b00000100100010011100001001001001;
12'b100000010100: dataA <= 32'b01010110101110100111101011010111;
12'b100000010101: dataA <= 32'b00000111000001100110001110000011;
12'b100000010110: dataA <= 32'b00000111100001000010110001101000;
12'b100000010111: dataA <= 32'b00001000010101101101010000111111;
12'b100000011000: dataA <= 32'b01111000011100110011101101101111;
12'b100000011001: dataA <= 32'b00000110101010100110100111010010;
12'b100000011010: dataA <= 32'b11011111000001110101100100110100;
12'b100000011011: dataA <= 32'b00000001111000110101101001010100;
12'b100000011100: dataA <= 32'b00110101010100110010000101100111;
12'b100000011101: dataA <= 32'b00000001001111010000111111100110;
12'b100000011110: dataA <= 32'b01110001000010101110101110011000;
12'b100000011111: dataA <= 32'b00000010011001010101011010010100;
12'b100000100000: dataA <= 32'b11110010010001010111100011011001;
12'b100000100001: dataA <= 32'b00000110000111100010001100011001;
12'b100000100010: dataA <= 32'b10010111000110101101010010110010;
12'b100000100011: dataA <= 32'b00001011000011100010001100101100;
12'b100000100100: dataA <= 32'b00011110011010101111010010110100;
12'b100000100101: dataA <= 32'b00001111010001010110110101010010;
12'b100000100110: dataA <= 32'b11110001001001001011100111001100;
12'b100000100111: dataA <= 32'b00000001101001001010010100100100;
12'b100000101000: dataA <= 32'b11010000001010110001110101000110;
12'b100000101001: dataA <= 32'b00000101111110100011101001100001;
12'b100000101010: dataA <= 32'b11101100100110000111100111010110;
12'b100000101011: dataA <= 32'b00001011000010110100010110001010;
12'b100000101100: dataA <= 32'b10010011000111001110110110010000;
12'b100000101101: dataA <= 32'b00000001101100100110110001111100;
12'b100000101110: dataA <= 32'b11001110111010100111101000011001;
12'b100000101111: dataA <= 32'b00001010100110001100010010011011;
12'b100000110000: dataA <= 32'b10000011000011001101100001010011;
12'b100000110001: dataA <= 32'b00000100110011101111001110010100;
12'b100000110010: dataA <= 32'b01111101001001010010111110001000;
12'b100000110011: dataA <= 32'b00000101110110001101010100111100;
12'b100000110100: dataA <= 32'b01011000010010010110011011110111;
12'b100000110101: dataA <= 32'b00001101001100110110011101100010;
12'b100000110110: dataA <= 32'b00111010100000100101000100110011;
12'b100000110111: dataA <= 32'b00001011010110011011001110111010;
12'b100000111000: dataA <= 32'b10000110100101000001110010000110;
12'b100000111001: dataA <= 32'b00000001010111001111011101110010;
12'b100000111010: dataA <= 32'b11010001101001100011101000101110;
12'b100000111011: dataA <= 32'b00001010001010010010001000101110;
12'b100000111100: dataA <= 32'b11101101000000011010011110101001;
12'b100000111101: dataA <= 32'b00001011010001100100111111110100;
12'b100000111110: dataA <= 32'b11010010101101101011001100101011;
12'b100000111111: dataA <= 32'b00000111110111101001011000001010;
12'b100001000000: dataA <= 32'b00011100110101011101111000010100;
12'b100001000001: dataA <= 32'b00001100111011000011000000010100;
12'b100001000010: dataA <= 32'b11101001011110001011110001101011;
12'b100001000011: dataA <= 32'b00000100010100011011001100101110;
12'b100001000100: dataA <= 32'b00110110100110001010010110001000;
12'b100001000101: dataA <= 32'b00000101000010101110001101000010;
12'b100001000110: dataA <= 32'b10000011000000111110000110010111;
12'b100001000111: dataA <= 32'b00001001100110011110010010111100;
12'b100001001000: dataA <= 32'b00010000111011110100000001101100;
12'b100001001001: dataA <= 32'b00000110000001001110001111000100;
12'b100001001010: dataA <= 32'b00101100110010000011000010000110;
12'b100001001011: dataA <= 32'b00000100101101111100110100110011;
12'b100001001100: dataA <= 32'b10010101011010100111101100111011;
12'b100001001101: dataA <= 32'b00001011010000111101000001100111;
12'b100001001110: dataA <= 32'b01101010100001000010010111001000;
12'b100001001111: dataA <= 32'b00001010101100011110101000111010;
12'b100001010000: dataA <= 32'b01001111010001110110011110011000;
12'b100001010001: dataA <= 32'b00000001001111110111000000110110;
12'b100001010010: dataA <= 32'b10000101000001001110010010010110;
12'b100001010011: dataA <= 32'b00000011111100000101010101001100;
12'b100001010100: dataA <= 32'b00100100110000010101101111010100;
12'b100001010101: dataA <= 32'b00000001010111000101001101101011;
12'b100001010110: dataA <= 32'b11100011001110001010101001000001;
12'b100001010111: dataA <= 32'b00001100100110001110010100111100;
12'b100001011000: dataA <= 32'b01101111011000110110101010011010;
12'b100001011001: dataA <= 32'b00001010101010110100101000010101;
12'b100001011010: dataA <= 32'b11100011010010011010000111000111;
12'b100001011011: dataA <= 32'b00001101010100010101000111001110;
12'b100001011100: dataA <= 32'b01001001001010110011011000001101;
12'b100001011101: dataA <= 32'b00001000010010010111000111110101;
12'b100001011110: dataA <= 32'b01011110111100011110000111110101;
12'b100001011111: dataA <= 32'b00000111000110101000001110011100;
12'b100001100000: dataA <= 32'b10010100111000110100101011010010;
12'b100001100001: dataA <= 32'b00000110011010101001100101111011;
12'b100001100010: dataA <= 32'b10100010001110100101000100110010;
12'b100001100011: dataA <= 32'b00001011111100101111010110101001;
12'b100001100100: dataA <= 32'b01010001100010010111101001010111;
12'b100001100101: dataA <= 32'b00000110011110011111011001101110;
12'b100001100110: dataA <= 32'b10100001010010010110100101010110;
12'b100001100111: dataA <= 32'b00001010001000110110100000001100;
12'b100001101000: dataA <= 32'b11010000001001100011000011101011;
12'b100001101001: dataA <= 32'b00000110000001100000001001011000;
12'b100001101010: dataA <= 32'b01011000101010001111101010011000;
12'b100001101011: dataA <= 32'b00001000100001101010010010000011;
12'b100001101100: dataA <= 32'b10000101010101001010010010100110;
12'b100001101101: dataA <= 32'b00000111110101101011010100101110;
12'b100001101110: dataA <= 32'b11111010100100110011001101110001;
12'b100001101111: dataA <= 32'b00000111001010101000101011011010;
12'b100001110000: dataA <= 32'b10011111000001101101100100010011;
12'b100001110001: dataA <= 32'b00000001010101101111101101010100;
12'b100001110010: dataA <= 32'b11110011011101000001100110100110;
12'b100001110011: dataA <= 32'b00000001101101010000110111010110;
12'b100001110100: dataA <= 32'b01110001001010011110111101011010;
12'b100001110101: dataA <= 32'b00000001110111010011010110010100;
12'b100001110110: dataA <= 32'b01110110011001000111000010010110;
12'b100001110111: dataA <= 32'b00000111000111100110001100101001;
12'b100001111000: dataA <= 32'b11010111000010100101100010101111;
12'b100001111001: dataA <= 32'b00001100000101100110001100101011;
12'b100001111010: dataA <= 32'b11100010011110010111100010010010;
12'b100001111011: dataA <= 32'b00001111010100010110110001100001;
12'b100001111100: dataA <= 32'b01110001010001001011010111001100;
12'b100001111101: dataA <= 32'b00000010100111001110001100100100;
12'b100001111110: dataA <= 32'b11010110000111000010010110000101;
12'b100001111111: dataA <= 32'b00000100011101011111101001110001;
12'b100010000000: dataA <= 32'b11101110101101101111100110110110;
12'b100010000001: dataA <= 32'b00001100000011111000011110010010;
12'b100010000010: dataA <= 32'b10010011000010111111010110010000;
12'b100010000011: dataA <= 32'b00000010001010101000110101111100;
12'b100010000100: dataA <= 32'b11001110110010001111100111011000;
12'b100010000101: dataA <= 32'b00001011100111010000001010011011;
12'b100010000110: dataA <= 32'b10000010110110111110000001010001;
12'b100010000111: dataA <= 32'b00000100110010101101010110010100;
12'b100010001000: dataA <= 32'b11111101010101011010101111001011;
12'b100010001001: dataA <= 32'b00000101010101001011001100111011;
12'b100010001010: dataA <= 32'b01011100010010000110011010111001;
12'b100010001011: dataA <= 32'b00001101101110111010100101101010;
12'b100010001100: dataA <= 32'b10111100101100011100100100110010;
12'b100010001101: dataA <= 32'b00001010010111011001001111001010;
12'b100010001110: dataA <= 32'b10001010011101010001100011000100;
12'b100010001111: dataA <= 32'b00000000110100001101010101111010;
12'b100010010000: dataA <= 32'b01001111100001100011011000101110;
12'b100010010001: dataA <= 32'b00001010101011011000000100100110;
12'b100010010010: dataA <= 32'b10101101001000101001111111001100;
12'b100010010011: dataA <= 32'b00001011010010100100111111101101;
12'b100010010100: dataA <= 32'b00010100101001110011001101001101;
12'b100010010101: dataA <= 32'b00000110110111100111011100010010;
12'b100010010110: dataA <= 32'b10011100110101001101100111110100;
12'b100010010111: dataA <= 32'b00001011111101000010110100010011;
12'b100010011000: dataA <= 32'b01100101100010001011110010001001;
12'b100010011001: dataA <= 32'b00000011110010011001001100100110;
12'b100010011010: dataA <= 32'b10111000101110010010010111001000;
12'b100010011011: dataA <= 32'b00000110100001110010010101010001;
12'b100010011100: dataA <= 32'b00000010110100101101100101010110;
12'b100010011101: dataA <= 32'b00001010100111100010010010111101;
12'b100010011110: dataA <= 32'b10010000110011110100110010001010;
12'b100010011111: dataA <= 32'b00000111100001010100001011000100;
12'b100010100000: dataA <= 32'b10101100110110001011000011000100;
12'b100010100001: dataA <= 32'b00000100101100111101000000111010;
12'b100010100010: dataA <= 32'b01010011010110001111101011111101;
12'b100010100011: dataA <= 32'b00001011010010111101001101001111;
12'b100010100100: dataA <= 32'b11101110100101010001111000001000;
12'b100010100101: dataA <= 32'b00001010101101100000101001001001;
12'b100010100110: dataA <= 32'b10001101001001100110011101011011;
12'b100010100111: dataA <= 32'b00000001101101110101001000100101;
12'b100010101000: dataA <= 32'b01000100111000111101110001110100;
12'b100010101001: dataA <= 32'b00000010011010000011001001001100;
12'b100010101010: dataA <= 32'b00100110110000001100111110110111;
12'b100010101011: dataA <= 32'b00000000110100000101000101110011;
12'b100010101100: dataA <= 32'b01100011001110010010101010100001;
12'b100010101101: dataA <= 32'b00001101101001010010001100111100;
12'b100010101110: dataA <= 32'b10101011100000101110001001011011;
12'b100010101111: dataA <= 32'b00001011001011110110110000001100;
12'b100010110000: dataA <= 32'b01100001010010101010011000000111;
12'b100010110001: dataA <= 32'b00001100110110010101000010111111;
12'b100010110010: dataA <= 32'b11001001000010110011101000001101;
12'b100010110011: dataA <= 32'b00001000010010010111000011100101;
12'b100010110100: dataA <= 32'b10011110111100010101010111010101;
12'b100010110101: dataA <= 32'b00001000000110101100010010011100;
12'b100010110110: dataA <= 32'b10010100110100110100001011010011;
12'b100010110111: dataA <= 32'b00000101011001100101101001111011;
12'b100010111000: dataA <= 32'b11100110001110011101010100110001;
12'b100010111001: dataA <= 32'b00001010011110101101011110111001;
12'b100010111010: dataA <= 32'b00001101011001111111101000010111;
12'b100010111011: dataA <= 32'b00000100111101011011011001011110;
12'b100010111100: dataA <= 32'b11011111010010000110100100110101;
12'b100010111101: dataA <= 32'b00001010101001111010101000001011;
12'b100010111110: dataA <= 32'b10010110000101101011000100001001;
12'b100010111111: dataA <= 32'b00000111100001100110001101110000;
12'b100011000000: dataA <= 32'b01011010101001110111101001011001;
12'b100011000001: dataA <= 32'b00001010000001101110010110001011;
12'b100011000010: dataA <= 32'b00000011001101010010000011100100;
12'b100011000011: dataA <= 32'b00000111010100101001011000011110;
12'b100011000100: dataA <= 32'b01111100110000111010101101010011;
12'b100011000101: dataA <= 32'b00000111101010101010101111100011;
12'b100011000110: dataA <= 32'b01011111000001011101010100010001;
12'b100011000111: dataA <= 32'b00000000110011101011110101001100;
12'b100011001000: dataA <= 32'b00101111100001010001010111100110;
12'b100011001001: dataA <= 32'b00000010001010010000110010111111;
12'b100011001010: dataA <= 32'b10101111010010001111001100011100;
12'b100011001011: dataA <= 32'b00000000110100010001001110010100;
12'b100011001100: dataA <= 32'b11111000100000101110100001110100;
12'b100011001101: dataA <= 32'b00001000000111101100010000111000;
12'b100011001110: dataA <= 32'b01010110111110010101110010101101;
12'b100011001111: dataA <= 32'b00001101000110101100010000101011;
12'b100011010000: dataA <= 32'b10100110011101111111100010010000;
12'b100011010001: dataA <= 32'b00001110110111011000101101110001;
12'b100011010010: dataA <= 32'b11101101011001010010110111101100;
12'b100011010011: dataA <= 32'b00000011000101010100001000011011;
12'b100011010100: dataA <= 32'b11011100000111001010100111000101;
12'b100011010101: dataA <= 32'b00000011011011011011100110000001;
12'b100011010110: dataA <= 32'b00110000110001010111100101110101;
12'b100011010111: dataA <= 32'b00001101000101111010101010011011;
12'b100011011000: dataA <= 32'b10010010111010100111100110001111;
12'b100011011001: dataA <= 32'b00000010101000101000110101110100;
12'b100011011010: dataA <= 32'b00010000101001110111100110011000;
12'b100011011011: dataA <= 32'b00001100101001010110000110011100;
12'b100011011100: dataA <= 32'b11000010101010101110100001001110;
12'b100011011101: dataA <= 32'b00000100010000101011011010001100;
12'b100011011110: dataA <= 32'b01111001011101100010011111001101;
12'b100011011111: dataA <= 32'b00000100110100001011000101000011;
12'b100011100000: dataA <= 32'b00100000001101110110011001111001;
12'b100011100001: dataA <= 32'b00001101110000111100110001111010;
12'b100011100010: dataA <= 32'b00111100111000011100000100010000;
12'b100011100011: dataA <= 32'b00001001111000011001001011001011;
12'b100011100100: dataA <= 32'b10001100010101100001010100100010;
12'b100011100101: dataA <= 32'b00000000110001001011001110000010;
12'b100011100110: dataA <= 32'b10001011011001100011011000101110;
12'b100011100111: dataA <= 32'b00001011001100011110000100010101;
12'b100011101000: dataA <= 32'b00101101001100110001011111001111;
12'b100011101001: dataA <= 32'b00001010110100100101000011100110;
12'b100011101010: dataA <= 32'b10010110100101110010111101001111;
12'b100011101011: dataA <= 32'b00000110010111100011011100100001;
12'b100011101100: dataA <= 32'b11011110110101000101010111010011;
12'b100011101101: dataA <= 32'b00001010011110000010101000011010;
12'b100011101110: dataA <= 32'b10100011100010001011110010100111;
12'b100011101111: dataA <= 32'b00000011110001011001001000010101;
12'b100011110000: dataA <= 32'b10111010111010100010100111100111;
12'b100011110001: dataA <= 32'b00001000000001110110011101100001;
12'b100011110010: dataA <= 32'b01000010101000100101000100110101;
12'b100011110011: dataA <= 32'b00001011101000100110010110110101;
12'b100011110100: dataA <= 32'b00010010101111101101100010101000;
12'b100011110101: dataA <= 32'b00001001000001011000000110111101;
12'b100011110110: dataA <= 32'b00101110111110001011000100100010;
12'b100011110111: dataA <= 32'b00000101001010111101001101000010;
12'b100011111000: dataA <= 32'b00010001001101110111101010011110;
12'b100011111001: dataA <= 32'b00001011010011111011011000111111;
12'b100011111010: dataA <= 32'b10110000101101011001101000101000;
12'b100011111011: dataA <= 32'b00001011001110100010101101010001;
12'b100011111100: dataA <= 32'b00001101000001010110001011111100;
12'b100011111101: dataA <= 32'b00000010001010110101010000011101;
12'b100011111110: dataA <= 32'b11000110101100101101010001010001;
12'b100011111111: dataA <= 32'b00000001110111000011000001001011;
12'b100100000000: dataA <= 32'b11100110110100001100001101111001;
12'b100100000001: dataA <= 32'b00000000110001000100111001110010;
12'b100100000010: dataA <= 32'b11100001001110011010111011100011;
12'b100100000011: dataA <= 32'b00001110001011010110001000111011;
12'b100100000100: dataA <= 32'b11101001100100011101011000011011;
12'b100100000101: dataA <= 32'b00001011101101111000111000001011;
12'b100100000110: dataA <= 32'b10011111010010110010101001001000;
12'b100100000111: dataA <= 32'b00001100010111010100111110100111;
12'b100100001000: dataA <= 32'b10001000111010110100001000101101;
12'b100100001001: dataA <= 32'b00000111110010010110111111010110;
12'b100100001010: dataA <= 32'b10011110111100001100110110110101;
12'b100100001011: dataA <= 32'b00001001000111110000010110011100;
12'b100100001100: dataA <= 32'b10010110110000110011101010110101;
12'b100100001101: dataA <= 32'b00000100111000100001101001111011;
12'b100100001110: dataA <= 32'b01101100010010010101010100101111;
12'b100100001111: dataA <= 32'b00001001011110101001100011001010;
12'b100100010000: dataA <= 32'b11001011010001100111100111110111;
12'b100100010001: dataA <= 32'b00000011111100011001011001001101;
12'b100100010010: dataA <= 32'b00011111010001110110100100010100;
12'b100100010011: dataA <= 32'b00001011001011111010110100001011;
12'b100100010100: dataA <= 32'b10011100000101110010110100101000;
12'b100100010101: dataA <= 32'b00001001000001101010010010000000;
12'b100100010110: dataA <= 32'b01011100100101011111101000011001;
12'b100100010111: dataA <= 32'b00001011100010110010011110001011;
12'b100100011000: dataA <= 32'b01000011000001100001110100100011;
12'b100100011001: dataA <= 32'b00000110110100100101011100010101;
12'b100100011010: dataA <= 32'b00111100111101000010001100110101;
12'b100100011011: dataA <= 32'b00001000001010101100110011100100;
12'b100100011100: dataA <= 32'b11011111000001010101000100010000;
12'b100100011101: dataA <= 32'b00000000110000100101110101001011;
12'b100100011110: dataA <= 32'b10101011101001100001001000100110;
12'b100100011111: dataA <= 32'b00000010101000010010101010101111;
12'b100100100000: dataA <= 32'b10101101010101111111001010111101;
12'b100100100001: dataA <= 32'b00000000110010001111001010001100;
12'b100100100010: dataA <= 32'b10111100101100011110000001010010;
12'b100100100011: dataA <= 32'b00001000100111110000010101010000;
12'b100100100100: dataA <= 32'b11010110111110001101110011001011;
12'b100100100101: dataA <= 32'b00001110001001110000010100110010;
12'b100100100110: dataA <= 32'b10101000100001101111100010001110;
12'b100100100111: dataA <= 32'b00001101111001011010101101111001;
12'b100100101000: dataA <= 32'b00101011011101011010101000001100;
12'b100100101001: dataA <= 32'b00000100100011011010000100100011;
12'b100100101010: dataA <= 32'b11100010000111010011001000100101;
12'b100100101011: dataA <= 32'b00000010011001010111100010001001;
12'b100100101100: dataA <= 32'b00110010111001000111000101010100;
12'b100100101101: dataA <= 32'b00001110001000111100110110011011;
12'b100100101110: dataA <= 32'b10010100110110001111100110101110;
12'b100100101111: dataA <= 32'b00000011100110101000111001110100;
12'b100100110000: dataA <= 32'b01010010100101011111100101110111;
12'b100100110001: dataA <= 32'b00001101001011011100000110010100;
12'b100100110010: dataA <= 32'b11000110100010011110100001001011;
12'b100100110011: dataA <= 32'b00000100001111101001011110001100;
12'b100100110100: dataA <= 32'b00110101101001101010011111010000;
12'b100100110101: dataA <= 32'b00000100010010001010111001000011;
12'b100100110110: dataA <= 32'b00100110010001100110001000111010;
12'b100100110111: dataA <= 32'b00001101010010111100111110000010;
12'b100100111000: dataA <= 32'b10111101000100011011010100001111;
12'b100100111001: dataA <= 32'b00001000111001010111000111010011;
12'b100100111010: dataA <= 32'b10010010001101110001000101100001;
12'b100100111011: dataA <= 32'b00000000101110001001000110001010;
12'b100100111100: dataA <= 32'b11001001010001101011001001001111;
12'b100100111101: dataA <= 32'b00001011001101100100000100001100;
12'b100100111110: dataA <= 32'b10101011010001001000111111010010;
12'b100100111111: dataA <= 32'b00001010010101100101000011010110;
12'b100101000000: dataA <= 32'b00011010100001111010111101010001;
12'b100101000001: dataA <= 32'b00000101010110100001011100110001;
12'b100101000010: dataA <= 32'b01011110110100111100110111010011;
12'b100101000011: dataA <= 32'b00001000111110000110100000100010;
12'b100101000100: dataA <= 32'b11011111100010001011110011100101;
12'b100101000101: dataA <= 32'b00000011101111010111000100001100;
12'b100101000110: dataA <= 32'b01111011000010101010111000101000;
12'b100101000111: dataA <= 32'b00001001000001111000100101110001;
12'b100101001000: dataA <= 32'b10000110100000100100010100010100;
12'b100101001001: dataA <= 32'b00001100001010101010011010100101;
12'b100101001010: dataA <= 32'b01010100101011100110000011100110;
12'b100101001011: dataA <= 32'b00001010100001011110000110110101;
12'b100101001100: dataA <= 32'b11101111000010010011000101100001;
12'b100101001101: dataA <= 32'b00000101101010111011011001010001;
12'b100101001110: dataA <= 32'b10001111001001011111101000111110;
12'b100101001111: dataA <= 32'b00001010110100111001100000101110;
12'b100101010000: dataA <= 32'b01110000110001101001101001001001;
12'b100101010001: dataA <= 32'b00001011010000100100101101100001;
12'b100101010010: dataA <= 32'b10001100111001000101111010111110;
12'b100101010011: dataA <= 32'b00000010101000110011011000010100;
12'b100101010100: dataA <= 32'b10001000100100101100110001001111;
12'b100101010101: dataA <= 32'b00000000110101000010110101001011;
12'b100101010110: dataA <= 32'b11101000111000001011011100111011;
12'b100101010111: dataA <= 32'b00000000101110000100101101111010;
12'b100101011000: dataA <= 32'b10011111001110100010111101000101;
12'b100101011001: dataA <= 32'b00001110101101011100000100111011;
12'b100101011010: dataA <= 32'b01100101100100010100110111011011;
12'b100101011011: dataA <= 32'b00001011101110111001000000001011;
12'b100101011100: dataA <= 32'b10011111010010111010111001101000;
12'b100101011101: dataA <= 32'b00001011011001010100111010001111;
12'b100101011110: dataA <= 32'b00001000110010110100011000101101;
12'b100101011111: dataA <= 32'b00000111110010010110111111000111;
12'b100101100000: dataA <= 32'b11011110111100001100000110010100;
12'b100101100001: dataA <= 32'b00001010000111110100011110010100;
12'b100101100010: dataA <= 32'b10010110101100111011001010010101;
12'b100101100011: dataA <= 32'b00000011110111011101101001111011;
12'b100101100100: dataA <= 32'b11110000010110001101100100101110;
12'b100101100101: dataA <= 32'b00000111111110100111100011010010;
12'b100101100110: dataA <= 32'b10001001001001001111010110110111;
12'b100101100111: dataA <= 32'b00000010111010010111010101000101;
12'b100101101000: dataA <= 32'b01011101010001100110010011110010;
12'b100101101001: dataA <= 32'b00001011101100111100111100010010;
12'b100101101010: dataA <= 32'b10100010000101111010110101100111;
12'b100101101011: dataA <= 32'b00001010100001110000010110011000;
12'b100101101100: dataA <= 32'b10011110100101000111010111111001;
12'b100101101101: dataA <= 32'b00001100100100110110100110010011;
12'b100101101110: dataA <= 32'b10000010110101110001110110000010;
12'b100101101111: dataA <= 32'b00000110010011100011011100001100;
12'b100101110000: dataA <= 32'b10111101001001010001111100010111;
12'b100101110001: dataA <= 32'b00001000101010101110110111100100;
12'b100101110010: dataA <= 32'b10011111000001001100110100001110;
12'b100101110011: dataA <= 32'b00000000101101100001111001001011;
12'b100101110100: dataA <= 32'b10100111101101111000111001100111;
12'b100101110101: dataA <= 32'b00000011000110010100100110010111;
12'b100101110110: dataA <= 32'b10101011011001100110111001011110;
12'b100101110111: dataA <= 32'b00000000101111001111000010001100;
12'b100101111000: dataA <= 32'b01111100110100010101100001001111;
12'b100101111001: dataA <= 32'b00001001100111110100011101101000;
12'b100101111010: dataA <= 32'b10010110111001111101110011101010;
12'b100101111011: dataA <= 32'b00001110101011110100011100111010;
12'b100101111100: dataA <= 32'b10101100100101010111010010101100;
12'b100101111101: dataA <= 32'b00001100111011011100101010001001;
12'b100101111110: dataA <= 32'b10101001100001100010011000101100;
12'b100101111111: dataA <= 32'b00000101100010100000000100101010;
12'b100110000000: dataA <= 32'b11101000000111010011101001100101;
12'b100110000001: dataA <= 32'b00000001010111010011011110011001;
12'b100110000010: dataA <= 32'b01110011000000101110100100110011;
12'b100110000011: dataA <= 32'b00001111001010111101000010100011;
12'b100110000100: dataA <= 32'b01010100110001110111100110101110;
12'b100110000101: dataA <= 32'b00000100100100101000111101101100;
12'b100110000110: dataA <= 32'b01010110100001000111010100110110;
12'b100110000111: dataA <= 32'b00001101001101100010000110010100;
12'b100110001000: dataA <= 32'b11001010010110001110110001101001;
12'b100110001001: dataA <= 32'b00000100101101100101100010000100;
12'b100110001010: dataA <= 32'b11110001110001111010001111010011;
12'b100110001011: dataA <= 32'b00000100010001001010110001001010;
12'b100110001100: dataA <= 32'b01101010010101010110000111111010;
12'b100110001101: dataA <= 32'b00001101010100111101001010010010;
12'b100110001110: dataA <= 32'b00111101010000100010110100101101;
12'b100110001111: dataA <= 32'b00000111111001010111000011010100;
12'b100110010000: dataA <= 32'b11010110001010001001000111000001;
12'b100110010001: dataA <= 32'b00000000101011001000111010010010;
12'b100110010010: dataA <= 32'b00000111001001110011001001001111;
12'b100110010011: dataA <= 32'b00001011101111101010000100001100;
12'b100110010100: dataA <= 32'b00101001010101011000101111010101;
12'b100110010101: dataA <= 32'b00001001110110100101000010111111;
12'b100110010110: dataA <= 32'b10011100100010000010111100110011;
12'b100110010111: dataA <= 32'b00000100110101011101011101000000;
12'b100110011000: dataA <= 32'b11100000110100111100010110110011;
12'b100110011001: dataA <= 32'b00000111011110001010010100110001;
12'b100110011010: dataA <= 32'b00011011100010001100000101000100;
12'b100110011011: dataA <= 32'b00000011101101010111000000001100;
12'b100110011100: dataA <= 32'b01111011001110110011001001001000;
12'b100110011101: dataA <= 32'b00001010100010111010110010000001;
12'b100110011110: dataA <= 32'b11001010010100011011110011110010;
12'b100110011111: dataA <= 32'b00001100101011101110011110011101;
12'b100110100000: dataA <= 32'b10010110100111010110100100100100;
12'b100110100001: dataA <= 32'b00001011100011100100000110101101;
12'b100110100010: dataA <= 32'b10101101001010011011010111000001;
12'b100110100011: dataA <= 32'b00000110101001111001100001011001;
12'b100110100100: dataA <= 32'b11001111000001000111010111011110;
12'b100110100101: dataA <= 32'b00001010010101110101101000011101;
12'b100110100110: dataA <= 32'b01110010111001111001101010001010;
12'b100110100111: dataA <= 32'b00001011010001100110110001110001;
12'b100110101000: dataA <= 32'b11001110110000111101011001011110;
12'b100110101001: dataA <= 32'b00000011000110101111011100010011;
12'b100110101010: dataA <= 32'b01001100011100100100010001001100;
12'b100110101011: dataA <= 32'b00000000110010000100101001001011;
12'b100110101100: dataA <= 32'b11101000111100001010111011111101;
12'b100110101101: dataA <= 32'b00000000101011000110100110000010;
12'b100110101110: dataA <= 32'b00011101001110101011001110000111;
12'b100110101111: dataA <= 32'b00001110110000100010000100111011;
12'b100110110000: dataA <= 32'b10100001100100010100000110011010;
12'b100110110001: dataA <= 32'b00001011110000110111001100010010;
12'b100110110010: dataA <= 32'b10011101010011000011011010001001;
12'b100110110011: dataA <= 32'b00001010011010010110110101110111;
12'b100110110100: dataA <= 32'b01001010101010110100101001001110;
12'b100110110101: dataA <= 32'b00000111110010010110111010110111;
12'b100110110110: dataA <= 32'b11011110111100001011010101110011;
12'b100110110111: dataA <= 32'b00001010101000110110101010001100;
12'b100110111000: dataA <= 32'b10011000101000111010101001010110;
12'b100110111001: dataA <= 32'b00000011010101011001100110000011;
12'b100110111010: dataA <= 32'b01110100011110000101100100101101;
12'b100110111011: dataA <= 32'b00000110011110100011100111010011;
12'b100110111100: dataA <= 32'b00001001000000111111000110010110;
12'b100110111101: dataA <= 32'b00000001110111010101010000111101;
12'b100110111110: dataA <= 32'b11011011001101010110000011110001;
12'b100110111111: dataA <= 32'b00001011101101111011001000011001;
12'b100111000000: dataA <= 32'b11101000000101111010110110100110;
12'b100111000001: dataA <= 32'b00001011100011110100011110101000;
12'b100111000010: dataA <= 32'b10100010100100110110110110111001;
12'b100111000011: dataA <= 32'b00001101100110111000101110010011;
12'b100111000100: dataA <= 32'b00000100101001111001110111100001;
12'b100111000101: dataA <= 32'b00000110010011011111100000001100;
12'b100111000110: dataA <= 32'b01111101010101100001101011011000;
12'b100111000111: dataA <= 32'b00001001001010101110111111011101;
12'b100111001000: dataA <= 32'b01011111000001001100100100001101;
12'b100111001001: dataA <= 32'b00000001001010011011110101010011;
12'b100111001010: dataA <= 32'b10100011101110001000111010000111;
12'b100111001011: dataA <= 32'b00000100000101011000100001111111;
12'b100111001100: dataA <= 32'b11101001011101010110101000011110;
12'b100111001101: dataA <= 32'b00000000101100001110111010000100;
12'b100111001110: dataA <= 32'b01111101000000001100110001001100;
12'b100111001111: dataA <= 32'b00001010101000110110100101111000;
12'b100111010000: dataA <= 32'b00011000110101110101110100001000;
12'b100111010001: dataA <= 32'b00001110101110110110100101000010;
12'b100111010010: dataA <= 32'b11101110101000111111000010101010;
12'b100111010011: dataA <= 32'b00001011111101011110101010011001;
12'b100111010100: dataA <= 32'b00100101100001101010011000101100;
12'b100111010101: dataA <= 32'b00000111000010100110000100110010;
12'b100111010110: dataA <= 32'b00101110001011010100011010100110;
12'b100111010111: dataA <= 32'b00000000110100010001011010101010;
12'b100111011000: dataA <= 32'b10110011000100011110000100110010;
12'b100111011001: dataA <= 32'b00001111001101111101001110100011;
12'b100111011010: dataA <= 32'b01010110101101011111100110101101;
12'b100111011011: dataA <= 32'b00000101100011101001000001101100;
12'b100111011100: dataA <= 32'b10011000011100110110110100010101;
12'b100111011101: dataA <= 32'b00001101101111101000000110010100;
12'b100111011110: dataA <= 32'b11001110001101111110110010100110;
12'b100111011111: dataA <= 32'b00000100101100100011100001111100;
12'b100111100000: dataA <= 32'b01101101110110000010001110110110;
12'b100111100001: dataA <= 32'b00000011101111001100101001010010;
12'b100111100010: dataA <= 32'b01101110011001001101100110111010;
12'b100111100011: dataA <= 32'b00001100110110111101010010011010;
12'b100111100100: dataA <= 32'b10111011011100101010010100101100;
12'b100111100101: dataA <= 32'b00000111011001010111000011010100;
12'b100111100110: dataA <= 32'b11011100001010011001011000100001;
12'b100111100111: dataA <= 32'b00000001001001001010110010011010;
12'b100111101000: dataA <= 32'b01000110111101110011001001001111;
12'b100111101001: dataA <= 32'b00001011110000101110001100001011;
12'b100111101010: dataA <= 32'b10100111011001110000101110010111;
12'b100111101011: dataA <= 32'b00001001010110100011000110101111;
12'b100111101100: dataA <= 32'b01100000011110001010111100010101;
12'b100111101101: dataA <= 32'b00000100010011011011011101011000;
12'b100111101110: dataA <= 32'b01100000110100111100000110010010;
12'b100111101111: dataA <= 32'b00000101111110001110001101000001;
12'b100111110000: dataA <= 32'b01011001011110001100000110000011;
12'b100111110001: dataA <= 32'b00000100001100010111000000001011;
12'b100111110010: dataA <= 32'b01111001010110110011011010001001;
12'b100111110011: dataA <= 32'b00001100000011111100111110010001;
12'b100111110100: dataA <= 32'b11001110001100100011010011110001;
12'b100111110101: dataA <= 32'b00001101001101110000100110010101;
12'b100111110110: dataA <= 32'b11011010100010111111000101100011;
12'b100111110111: dataA <= 32'b00001101000101101010001010100101;
12'b100111111000: dataA <= 32'b01101101001110011011101000100001;
12'b100111111001: dataA <= 32'b00000111001000110101101001101001;
12'b100111111010: dataA <= 32'b01001110111000110110110101111110;
12'b100111111011: dataA <= 32'b00001001110110101111110000001101;
12'b100111111100: dataA <= 32'b01110011000010001001101010101010;
12'b100111111101: dataA <= 32'b00001010110010100110110010001001;
12'b100111111110: dataA <= 32'b00001110101100110100110111111110;
12'b100111111111: dataA <= 32'b00000100000101101101100100010011;
12'b101000000000: dataA <= 32'b00010000010100100011110001101010;
12'b101000000001: dataA <= 32'b00000000101111000110011101010011;
12'b101000000010: dataA <= 32'b11101000111100011010001010011110;
12'b101000000011: dataA <= 32'b00000001001000001010011010001010;
12'b101000000100: dataA <= 32'b10011101001110101011101110101001;
12'b101000000101: dataA <= 32'b00001110110011101000001001000010;
12'b101000000110: dataA <= 32'b11011101100100010011100101011010;
12'b101000000111: dataA <= 32'b00001011110001110101010100011001;
12'b101000001000: dataA <= 32'b10011011001111000011101011001010;
12'b101000001001: dataA <= 32'b00001001011011010110110001011111;
12'b101000001010: dataA <= 32'b10001110100010101100111001001110;
12'b101000001011: dataA <= 32'b00000111010001011000110110011111;
12'b101000001100: dataA <= 32'b11011110111100010010100101010010;
12'b101000001101: dataA <= 32'b00001011001001111000110010001100;
12'b101000001110: dataA <= 32'b10011100101001001010011000110111;
12'b101000001111: dataA <= 32'b00000010110011010101100010000011;
12'b101000010000: dataA <= 32'b11110110100101110101100101001100;
12'b101000010001: dataA <= 32'b00000100111101011111100111011011;
12'b101000010010: dataA <= 32'b10001000111000101110100101110101;
12'b101000010011: dataA <= 32'b00000000110101010011001100110100;
12'b101000010100: dataA <= 32'b00011001001101000101110011101111;
12'b101000010101: dataA <= 32'b00001100001111111011010100101001;
12'b101000010110: dataA <= 32'b01101110001010000010110111100101;
12'b101000010111: dataA <= 32'b00001101000100110110100111000001;
12'b101000011000: dataA <= 32'b11100100101000100110010101111000;
12'b101000011001: dataA <= 32'b00001110101000111010111010010011;
12'b101000011010: dataA <= 32'b01000110011110001001111000100001;
12'b101000011011: dataA <= 32'b00000101110010011101011100001011;
12'b101000011100: dataA <= 32'b11111001011101110001101010111001;
12'b101000011101: dataA <= 32'b00001001101011101111000011010101;
12'b101000011110: dataA <= 32'b00011111000001001100010100101011;
12'b101000011111: dataA <= 32'b00000001100111010101110101010011;
12'b101000100000: dataA <= 32'b10011111101110011001001011001000;
12'b101000100001: dataA <= 32'b00000101100011011010100001100111;
12'b101000100010: dataA <= 32'b11100101100001000110010110111110;
12'b101000100011: dataA <= 32'b00000001001001001110110101111100;
12'b101000100100: dataA <= 32'b01111101001100001100000001101010;
12'b101000100101: dataA <= 32'b00001011001001111000110010010000;
12'b101000100110: dataA <= 32'b11011000110001100101110101000111;
12'b101000100111: dataA <= 32'b00001110110001111000110001010001;
12'b101000101000: dataA <= 32'b00110000110000101110100011101000;
12'b101000101001: dataA <= 32'b00001010011110100000101010100010;
12'b101000101010: dataA <= 32'b10100001100101110010011001001101;
12'b101000101011: dataA <= 32'b00001000100010101010001001000001;
12'b101000101100: dataA <= 32'b01110010010011010100111011000111;
12'b101000101101: dataA <= 32'b00000000110001001111010010110010;
12'b101000101110: dataA <= 32'b11110001001100010101100100110001;
12'b101000101111: dataA <= 32'b00001111010000111011010110101011;
12'b101000110000: dataA <= 32'b00011000101001000111010111001101;
12'b101000110001: dataA <= 32'b00000111000010101001000101101100;
12'b101000110010: dataA <= 32'b10011100011100100110010011110011;
12'b101000110011: dataA <= 32'b00001101110001101110001010001100;
12'b101000110100: dataA <= 32'b11010010001001101110110011100101;
12'b101000110101: dataA <= 32'b00000101001011011111100001110100;
12'b101000110110: dataA <= 32'b00100111111010010010011101111001;
12'b101000110111: dataA <= 32'b00000100001110001110100101011010;
12'b101000111000: dataA <= 32'b10110010100001000101010101111001;
12'b101000111001: dataA <= 32'b00001011111000111001011110100010;
12'b101000111010: dataA <= 32'b00110111100100111001110101001011;
12'b101000111011: dataA <= 32'b00000110011000010110111111001101;
12'b101000111100: dataA <= 32'b00100010001010101001101010000001;
12'b101000111101: dataA <= 32'b00000010000110001100101010100011;
12'b101000111110: dataA <= 32'b11000110110101111010111001010000;
12'b101000111111: dataA <= 32'b00001011010010110100010000001010;
12'b101001000000: dataA <= 32'b10100101011010001000101101111010;
12'b101001000001: dataA <= 32'b00001000110110100011000110010111;
12'b101001000010: dataA <= 32'b01100010100010001011001011110111;
12'b101001000011: dataA <= 32'b00000100010010010111011001110000;
12'b101001000100: dataA <= 32'b00100010110100111011100110010010;
12'b101001000101: dataA <= 32'b00000100011101010010001001010001;
12'b101001000110: dataA <= 32'b11010101011010001100000111100010;
12'b101001000111: dataA <= 32'b00000100101010010110111100001010;
12'b101001001000: dataA <= 32'b10110101100010110011101010101010;
12'b101001001001: dataA <= 32'b00001101000101111101000110100001;
12'b101001001010: dataA <= 32'b00010010001000101010100011101111;
12'b101001001011: dataA <= 32'b00001101001111110010101010000110;
12'b101001001100: dataA <= 32'b00011100100010101111100111000010;
12'b101001001101: dataA <= 32'b00001110000111110000001110010110;
12'b101001001110: dataA <= 32'b01101011010010011011101010000001;
12'b101001001111: dataA <= 32'b00000111101000101111110001111001;
12'b101001010000: dataA <= 32'b10001110110100100110010100011101;
12'b101001010001: dataA <= 32'b00001001010110101011111000001100;
12'b101001010010: dataA <= 32'b01110011001010011001101011001100;
12'b101001010011: dataA <= 32'b00001010110011101000110110011001;
12'b101001010100: dataA <= 32'b10010000100100110100010110011110;
12'b101001010101: dataA <= 32'b00000101100011101001101000011010;
12'b101001010110: dataA <= 32'b11010100010000100011010010100111;
12'b101001010111: dataA <= 32'b00000000101100001010010101011010;
12'b101001011000: dataA <= 32'b00101001000000100001101000111110;
12'b101001011001: dataA <= 32'b00000010000110001110010110001011;
12'b101001011010: dataA <= 32'b01011011001010110011111111001100;
12'b101001011011: dataA <= 32'b00001110010101101100001101001010;
12'b101001011100: dataA <= 32'b01011001100100011010110100011000;
12'b101001011101: dataA <= 32'b00001011110011110011011100101001;
12'b101001011110: dataA <= 32'b01011001001111000100001011101011;
12'b101001011111: dataA <= 32'b00001000011011011000101101000111;
12'b101001100000: dataA <= 32'b10010000011010100101001001001111;
12'b101001100001: dataA <= 32'b00000111010001011000110010000111;
12'b101001100010: dataA <= 32'b00011110111100011001110101010001;
12'b101001100011: dataA <= 32'b00001100001011111010111110000101;
12'b101001100100: dataA <= 32'b10011110100101010010001000010111;
12'b101001100101: dataA <= 32'b00000010010001010001011110000011;
12'b101001100110: dataA <= 32'b01111000110001101101010101101011;
12'b101001100111: dataA <= 32'b00000011011011011011100111011100;
12'b101001101000: dataA <= 32'b00001010101100011101110101010100;
12'b101001101001: dataA <= 32'b00000000110010010011001000101100;
12'b101001101010: dataA <= 32'b11011001001000111101010011101101;
12'b101001101011: dataA <= 32'b00001100010001110111011101000000;
12'b101001101100: dataA <= 32'b10110010010010001010111000100101;
12'b101001101101: dataA <= 32'b00001110000111111000101111010001;
12'b101001101110: dataA <= 32'b11100110101000010101100100110111;
12'b101001101111: dataA <= 32'b00001111001011111011000010010011;
12'b101001110000: dataA <= 32'b10001010010110011001111010000010;
12'b101001110001: dataA <= 32'b00000101110001011001011100010010;
12'b101001110010: dataA <= 32'b01110101101010000001011001111010;
12'b101001110011: dataA <= 32'b00001010001100101111001011000110;
12'b101001110100: dataA <= 32'b11011111000001000011110101001010;
12'b101001110101: dataA <= 32'b00000010100101010001101101011010;
12'b101001110110: dataA <= 32'b01011011101110101001011011101010;
12'b101001110111: dataA <= 32'b00000110100011011110100001001111;
12'b101001111000: dataA <= 32'b11100001100000110101110101011101;
12'b101001111001: dataA <= 32'b00000010000111010000101101111100;
12'b101001111010: dataA <= 32'b10111011011000001011010010101000;
12'b101001111011: dataA <= 32'b00001011101011111000111010101000;
12'b101001111100: dataA <= 32'b10011010110001011101100110000110;
12'b101001111101: dataA <= 32'b00001110110011111000111001100001;
12'b101001111110: dataA <= 32'b01110000111000011110000100100110;
12'b101001111111: dataA <= 32'b00001000111110100010101010110010;
12'b101010000000: dataA <= 32'b01011101100110000010001001001101;
12'b101010000001: dataA <= 32'b00001001100010110000001101001001;
12'b101010000010: dataA <= 32'b11110110011011001101011100001001;
12'b101010000011: dataA <= 32'b00000000101110001101001010111010;
12'b101010000100: dataA <= 32'b00101111010100001100110100001111;
12'b101010000101: dataA <= 32'b00001111010011111001100010101100;
12'b101010000110: dataA <= 32'b00011010101000110110110111001101;
12'b101010000111: dataA <= 32'b00001000000010101001001001101100;
12'b101010001000: dataA <= 32'b10100000011000010101100011110001;
12'b101010001001: dataA <= 32'b00001101010011110010010010001100;
12'b101010001010: dataA <= 32'b11011000000101011110100100100011;
12'b101010001011: dataA <= 32'b00000101101010011011100001110100;
12'b101010001100: dataA <= 32'b00100001111010011010011101011011;
12'b101010001101: dataA <= 32'b00000100001100010010011101101010;
12'b101010001110: dataA <= 32'b11110100100100111100110100111000;
12'b101010001111: dataA <= 32'b00001010111001110111100110101010;
12'b101010010000: dataA <= 32'b10110011101101000001010101101010;
12'b101010010001: dataA <= 32'b00000101010111010110111011000101;
12'b101010010010: dataA <= 32'b01100110001010111001111011100010;
12'b101010010011: dataA <= 32'b00000011000100001110100010100011;
12'b101010010100: dataA <= 32'b00001000101110000010111001010000;
12'b101010010101: dataA <= 32'b00001011010011111000011100011010;
12'b101010010110: dataA <= 32'b10100001011010011000101100011100;
12'b101010010111: dataA <= 32'b00000111110111100011000101111111;
12'b101010011000: dataA <= 32'b01100110100010010011001010111000;
12'b101010011001: dataA <= 32'b00000100010000010101010110001000;
12'b101010011010: dataA <= 32'b11100010110100111011000110010001;
12'b101010011011: dataA <= 32'b00000011011011011000000101100000;
12'b101010011100: dataA <= 32'b00010011010110001100001000100010;
12'b101010011101: dataA <= 32'b00000101001001010110111000011010;
12'b101010011110: dataA <= 32'b11110011101010111100001011001011;
12'b101010011111: dataA <= 32'b00001110000111111011010010110001;
12'b101010100000: dataA <= 32'b00011000000100110010000011101101;
12'b101010100001: dataA <= 32'b00001101010010110100110001110110;
12'b101010100010: dataA <= 32'b00100000011110010111101000000010;
12'b101010100011: dataA <= 32'b00001110101001110100010110000110;
12'b101010100100: dataA <= 32'b01101001010110011011111011100010;
12'b101010100101: dataA <= 32'b00001000101000101011111010010001;
12'b101010100110: dataA <= 32'b11010000101100010101100011011011;
12'b101010100111: dataA <= 32'b00001000010110100101111000001011;
12'b101010101000: dataA <= 32'b10110001010010101001111011001101;
12'b101010101001: dataA <= 32'b00001010010100101000111010101001;
12'b101010101010: dataA <= 32'b00010100100000101011110100111101;
12'b101010101011: dataA <= 32'b00000110100011100101101000101010;
12'b101010101100: dataA <= 32'b10011000001100101010110011000101;
12'b101010101101: dataA <= 32'b00000001001001001110001101100010;
12'b101010101110: dataA <= 32'b00101001000100110001000111011110;
12'b101010101111: dataA <= 32'b00000011000100010010001110010011;
12'b101010110000: dataA <= 32'b00011011001010110100001111001111;
12'b101010110001: dataA <= 32'b00001101010111110000010101011010;
12'b101010110010: dataA <= 32'b11010101100000100010010011010110;
12'b101010110011: dataA <= 32'b00001011010100101111100100111000;
12'b101010110100: dataA <= 32'b11011001001011000100101011101101;
12'b101010110101: dataA <= 32'b00000111011011011010101100110110;
12'b101010110110: dataA <= 32'b10010100010110011101011001001111;
12'b101010110111: dataA <= 32'b00000111010001011010110001101111;
12'b101010111000: dataA <= 32'b00011110111100101001010101010000;
12'b101010111001: dataA <= 32'b00001100001101111011000101111101;
12'b101010111010: dataA <= 32'b10100000100101100001110111010111;
12'b101010111011: dataA <= 32'b00000010001111001111010110000011;
12'b101010111100: dataA <= 32'b11111000111001100101010110001010;
12'b101010111101: dataA <= 32'b00000010011010010111100011010100;
12'b101010111110: dataA <= 32'b10001100100100001101010100110011;
12'b101010111111: dataA <= 32'b00000000101111010011000000101011;
endcase
if (enB)
case(addrB)
12'b000000000000: dataB <= 32'b11100101001110101110000110111000;
12'b000000000001: dataB <= 32'b00001000100111101110010000011101;
12'b000000000010: dataB <= 32'b01001000011001011011100010101110;
12'b000000000011: dataB <= 32'b00000011100011010110001100110001;
12'b000000000100: dataB <= 32'b01010100110010110111011011110110;
12'b000000000101: dataB <= 32'b00000101100001100000001001111011;
12'b000000000110: dataB <= 32'b01001011101000111011000001001011;
12'b000000000111: dataB <= 32'b00001000110100101111001101010111;
12'b000000001000: dataB <= 32'b11110100010100101011111101001100;
12'b000000001001: dataB <= 32'b00000110001011100100100011001001;
12'b000000001010: dataB <= 32'b00100001000001111101110101010101;
12'b000000001011: dataB <= 32'b00000010111010110111011101011101;
12'b000000001100: dataB <= 32'b10110111001000101010100101001000;
12'b000000001101: dataB <= 32'b00000001110010010001000011101101;
12'b000000001110: dataB <= 32'b00110000111110111110011110110101;
12'b000000001111: dataB <= 32'b00000011111011010111011110011100;
12'b000000010000: dataB <= 32'b10101100001001101111100100011010;
12'b000000010001: dataB <= 32'b00000101101000011100001100010010;
12'b000000010010: dataB <= 32'b11011001001010110101000011010011;
12'b000000010011: dataB <= 32'b00001001100010011100001100110100;
12'b000000010100: dataB <= 32'b01011100011111000111000011010110;
12'b000000010101: dataB <= 32'b00001111001110010100111001001010;
12'b000000010110: dataB <= 32'b10110011000101000011110110101101;
12'b000000010111: dataB <= 32'b00000001001100000110011100101101;
12'b000000011000: dataB <= 32'b00001100010010101001100100100111;
12'b000000011001: dataB <= 32'b00000111011110100101100101011010;
12'b000000011010: dataB <= 32'b10101010100010011111100111110111;
12'b000000011011: dataB <= 32'b00001001100001110000001110000010;
12'b000000011100: dataB <= 32'b10010101001011011110010110110001;
12'b000000011101: dataB <= 32'b00000001001111100100101110000100;
12'b000000011110: dataB <= 32'b10001100111110110111011000111000;
12'b000000011111: dataB <= 32'b00001001100101001000011010010011;
12'b000000100000: dataB <= 32'b01000011001111010101000001110110;
12'b000000100001: dataB <= 32'b00000101010100110001001010011100;
12'b000000100010: dataB <= 32'b10111100111101001011001101100101;
12'b000000100011: dataB <= 32'b00000110010111001111011001000100;
12'b000000100100: dataB <= 32'b10010010010110011110001100010110;
12'b000000100101: dataB <= 32'b00001100101010110010010001011010;
12'b000000100110: dataB <= 32'b11110110011000101101110101010100;
12'b000000100111: dataB <= 32'b00001011110101011101010010110001;
12'b000000101000: dataB <= 32'b11000100110000111010000001001000;
12'b000000101001: dataB <= 32'b00000010011001010001100001101010;
12'b000000101010: dataB <= 32'b00010111101101011011111000001101;
12'b000000101011: dataB <= 32'b00001001101001001110001101000111;
12'b000000101100: dataB <= 32'b00101100111100010011001110000111;
12'b000000101101: dataB <= 32'b00001011110000100010111011110100;
12'b000000101110: dataB <= 32'b10010000110001100011011100001010;
12'b000000101111: dataB <= 32'b00001000010111101011010100001011;
12'b000000110000: dataB <= 32'b11011010111001100110001000110011;
12'b000000110001: dataB <= 32'b00001101111001000011001100011100;
12'b000000110010: dataB <= 32'b00101011011010000011100001001110;
12'b000000110011: dataB <= 32'b00000100110101011101010001000111;
12'b000000110100: dataB <= 32'b01110100011010000010000101101001;
12'b000000110101: dataB <= 32'b00000011100011101000001000111010;
12'b000000110110: dataB <= 32'b01000011001101000110010110111000;
12'b000000110111: dataB <= 32'b00001001000101011000010111000100;
12'b000000111000: dataB <= 32'b11001110111111110011010001001111;
12'b000000111001: dataB <= 32'b00000100100010001010010111000011;
12'b000000111010: dataB <= 32'b01101010101101111011000001001000;
12'b000000111011: dataB <= 32'b00000100001110111100101000101011;
12'b000000111100: dataB <= 32'b10010111011110110111011101111001;
12'b000000111101: dataB <= 32'b00001011001111111100110101111111;
12'b000000111110: dataB <= 32'b10101000011100111010100110101001;
12'b000000111111: dataB <= 32'b00001010001011011100101100110010;
12'b000001000000: dataB <= 32'b10010001010101111110101110110110;
12'b000001000001: dataB <= 32'b00000001110010110100110101000110;
12'b000001000010: dataB <= 32'b11000111001101011110100010111001;
12'b000001000011: dataB <= 32'b00000100111101000111100001010100;
12'b000001000100: dataB <= 32'b01100010101100100110011111010001;
12'b000001000101: dataB <= 32'b00000010011001000111011001100011;
12'b000001000110: dataB <= 32'b00100101001010000010010111100001;
12'b000001000111: dataB <= 32'b00001011100101001010011101000101;
12'b000001001000: dataB <= 32'b00110001010101001110111011011001;
12'b000001001001: dataB <= 32'b00001010001001110010100000011110;
12'b000001001010: dataB <= 32'b01100101001110010001110110101000;
12'b000001001011: dataB <= 32'b00001101110001010111001011011110;
12'b000001001100: dataB <= 32'b10001011010110101011000111101101;
12'b000001001101: dataB <= 32'b00001000110001011001001011110100;
12'b000001001110: dataB <= 32'b00011111000000101110101000010101;
12'b000001001111: dataB <= 32'b00000110100111100010001010100100;
12'b000001010000: dataB <= 32'b11010010111100111100111011110001;
12'b000001010001: dataB <= 32'b00000111111011101011100001110011;
12'b000001010010: dataB <= 32'b01011100001110101100110101010011;
12'b000001010011: dataB <= 32'b00001101011011110001010010011001;
12'b000001010100: dataB <= 32'b10010011100110101111101001110110;
12'b000001010101: dataB <= 32'b00000111111110100001011001110110;
12'b000001010110: dataB <= 32'b10100111001110111101110111111000;
12'b000001010111: dataB <= 32'b00000111100111101010001000100110;
12'b000001011000: dataB <= 32'b11000100100001011011110010110000;
12'b000001011001: dataB <= 32'b00000010000101010010010000101001;
12'b000001011010: dataB <= 32'b01010100110111001110111100010100;
12'b000001011011: dataB <= 32'b00000100000010011100001001111011;
12'b000001011100: dataB <= 32'b10001111110000111011100000101110;
12'b000001011101: dataB <= 32'b00001001010100101111000101101111;
12'b000001011110: dataB <= 32'b01101110001100110100011100101010;
12'b000001011111: dataB <= 32'b00000101101100100000100010111001;
12'b000001100000: dataB <= 32'b01100001000010001101100101110110;
12'b000001100001: dataB <= 32'b00000011111100111011010101100101;
12'b000001100010: dataB <= 32'b11110111000000100011000100001001;
12'b000001100011: dataB <= 32'b00000001110100010001001011110100;
12'b000001100100: dataB <= 32'b00110000110111001101111111010010;
12'b000001100101: dataB <= 32'b00000100111101011011100010011100;
12'b000001100110: dataB <= 32'b01100110000110000111100101011100;
12'b000001100111: dataB <= 32'b00000100101001011000001100001011;
12'b000001101000: dataB <= 32'b01011001001110111100110011110101;
12'b000001101001: dataB <= 32'b00001000100010011000001100111101;
12'b000001101010: dataB <= 32'b11011000011111010110100100011000;
12'b000001101011: dataB <= 32'b00001111001011010100111101000010;
12'b000001101100: dataB <= 32'b11110010111101001100010110101101;
12'b000001101101: dataB <= 32'b00000001001110000100101000110101;
12'b000001101110: dataB <= 32'b01001000011010011001010011101001;
12'b000001101111: dataB <= 32'b00001000111110101001100001001010;
12'b000001110000: dataB <= 32'b10100110011110110111011000110110;
12'b000001110001: dataB <= 32'b00001000000001101010001001111010;
12'b000001110010: dataB <= 32'b10010101001111101101110110110001;
12'b000001110011: dataB <= 32'b00000001010001100010101110000100;
12'b000001110100: dataB <= 32'b10001111000111001110111001111000;
12'b000001110101: dataB <= 32'b00001000100100000100100010010011;
12'b000001110110: dataB <= 32'b01000101011011011100100010111000;
12'b000001110111: dataB <= 32'b00000101110101110001000010011100;
12'b000001111000: dataB <= 32'b00111100110001001011011100100100;
12'b000001111001: dataB <= 32'b00000111010111010011100001000101;
12'b000001111010: dataB <= 32'b11010000011010101101111100110100;
12'b000001111011: dataB <= 32'b00001100001000101110001101010010;
12'b000001111100: dataB <= 32'b10110010010000111110000101110101;
12'b000001111101: dataB <= 32'b00001100010011011111010010100001;
12'b000001111110: dataB <= 32'b11000100111000110010100000101011;
12'b000001111111: dataB <= 32'b00000011011011010101100101100010;
12'b000010000000: dataB <= 32'b10011011110001011100001000001101;
12'b000010000001: dataB <= 32'b00001001001001001000010101011111;
12'b000010000010: dataB <= 32'b01101100110100010011101101000100;
12'b000010000011: dataB <= 32'b00001011001110100010111011110011;
12'b000010000100: dataB <= 32'b01010000111001100011101011101000;
12'b000010000101: dataB <= 32'b00001001010111101101010000001100;
12'b000010000110: dataB <= 32'b01011010111001110110001001010011;
12'b000010000111: dataB <= 32'b00001110110111000101011000100101;
12'b000010001000: dataB <= 32'b10101101010110000011100001010000;
12'b000010001001: dataB <= 32'b00000101010110011111010001011111;
12'b000010001010: dataB <= 32'b11110000010101110010010101001010;
12'b000010001011: dataB <= 32'b00000010100101100010000100110010;
12'b000010001100: dataB <= 32'b11000101011001010110100111111000;
12'b000010001101: dataB <= 32'b00000111100101010100011011000011;
12'b000010001110: dataB <= 32'b01010001000111110010100001010001;
12'b000010001111: dataB <= 32'b00000011100011000110011111000011;
12'b000010010000: dataB <= 32'b00101000101001110011000000101011;
12'b000010010001: dataB <= 32'b00000100010000111000100000101100;
12'b000010010010: dataB <= 32'b10011011100011001110111110110111;
12'b000010010011: dataB <= 32'b00001011001101111100101010010111;
12'b000010010100: dataB <= 32'b00100100011000110011000110001001;
12'b000010010101: dataB <= 32'b00001001101010011010101100101011;
12'b000010010110: dataB <= 32'b00010011011110001110011111010011;
12'b000010010111: dataB <= 32'b00000001110100110100101101010111;
12'b000010011000: dataB <= 32'b00001001010101101110110011111010;
12'b000010011001: dataB <= 32'b00000110011110001011101001011101;
12'b000010011010: dataB <= 32'b10100000101100110110111111001110;
12'b000010011011: dataB <= 32'b00000011011011001011100001100011;
12'b000010011100: dataB <= 32'b10100101001001111010010110000001;
12'b000010011101: dataB <= 32'b00001010100011000110100101001101;
12'b000010011110: dataB <= 32'b10110011001101011111001100010111;
12'b000010011111: dataB <= 32'b00001001101000101110011000101110;
12'b000010100000: dataB <= 32'b11100111001110000001110101101000;
12'b000010100001: dataB <= 32'b00001101101111010111001111101101;
12'b000010100010: dataB <= 32'b11001101011110100010110111101101;
12'b000010100011: dataB <= 32'b00001000110001011001001111110011;
12'b000010100100: dataB <= 32'b11011111000000111111001000110101;
12'b000010100101: dataB <= 32'b00000101100111011110001010100011;
12'b000010100110: dataB <= 32'b11010011000001000101011011101111;
12'b000010100111: dataB <= 32'b00001000111011101111011101110011;
12'b000010101000: dataB <= 32'b00011000001110101100100101110100;
12'b000010101001: dataB <= 32'b00001101111001110011001010001001;
12'b000010101010: dataB <= 32'b10010111101010111111001010010101;
12'b000010101011: dataB <= 32'b00001001011110100101011010000110;
12'b000010101100: dataB <= 32'b00100111001011000101011000111000;
12'b000010101101: dataB <= 32'b00000110101000100100001000111111;
12'b000010101110: dataB <= 32'b10000010101101011100000011010010;
12'b000010101111: dataB <= 32'b00000001101000001110010100011010;
12'b000010110000: dataB <= 32'b01010010111011011110011100110010;
12'b000010110001: dataB <= 32'b00000011000100010110001101110011;
12'b000010110010: dataB <= 32'b10010101110100111100000000110000;
12'b000010110011: dataB <= 32'b00001001110011110001000010000111;
12'b000010110100: dataB <= 32'b00101010000100110100111100001001;
12'b000010110101: dataB <= 32'b00000101001101011110100010101001;
12'b000010110110: dataB <= 32'b01100001000010010101100110110111;
12'b000010110111: dataB <= 32'b00000101011101111011001001101101;
12'b000010111000: dataB <= 32'b00110110111000011011100011101011;
12'b000010111001: dataB <= 32'b00000010110111010001001111110100;
12'b000010111010: dataB <= 32'b11101110101111010101011111001111;
12'b000010111011: dataB <= 32'b00000110011110011101100010011011;
12'b000010111100: dataB <= 32'b00100000000110011111100110011101;
12'b000010111101: dataB <= 32'b00000100001010010010010000001100;
12'b000010111110: dataB <= 32'b11011011001110111100010100010111;
12'b000010111111: dataB <= 32'b00000111000010010010010001000101;
12'b000011000000: dataB <= 32'b00010100100011100110000101011010;
12'b000011000001: dataB <= 32'b00001110101000010101000000111011;
12'b000011000010: dataB <= 32'b01110000110101001100100110001110;
12'b000011000011: dataB <= 32'b00000001010001000010110001000110;
12'b000011000100: dataB <= 32'b10000100100010001001010011001010;
12'b000011000101: dataB <= 32'b00001010011110101101011101000010;
12'b000011000110: dataB <= 32'b11100010011011000111001001010110;
12'b000011000111: dataB <= 32'b00000110100001100110000101110010;
12'b000011001000: dataB <= 32'b10010111010011110101000110110010;
12'b000011001001: dataB <= 32'b00000001110100100000101110001100;
12'b000011001010: dataB <= 32'b01001111001111011110011010110111;
12'b000011001011: dataB <= 32'b00000111100100000010101110010011;
12'b000011001100: dataB <= 32'b00000111100011011100000011011010;
12'b000011001101: dataB <= 32'b00000110010110110000111010011100;
12'b000011001110: dataB <= 32'b01111010100101000011111011000010;
12'b000011001111: dataB <= 32'b00000111111000010101100101001101;
12'b000011010000: dataB <= 32'b00001100100010110101101101010010;
12'b000011010001: dataB <= 32'b00001011000110101000000101001011;
12'b000011010010: dataB <= 32'b01101110001001001110100110010110;
12'b000011010011: dataB <= 32'b00001100110001100001010010010001;
12'b000011010100: dataB <= 32'b00000101000100101011000000101110;
12'b000011010101: dataB <= 32'b00000100111101011001101001011011;
12'b000011010110: dataB <= 32'b10011111110001100100010111101101;
12'b000011010111: dataB <= 32'b00001000001000000110100001101111;
12'b000011011000: dataB <= 32'b10101100110000010100011011100011;
12'b000011011001: dataB <= 32'b00001011001101100010111011110010;
12'b000011011010: dataB <= 32'b00001110111101011011101010100111;
12'b000011011011: dataB <= 32'b00001001110111101111001000001101;
12'b000011011100: dataB <= 32'b11011010111110000110001001010011;
12'b000011011101: dataB <= 32'b00001111010100000111100000101101;
12'b000011011110: dataB <= 32'b10101111001110000011100001110011;
12'b000011011111: dataB <= 32'b00000110010111100001010001101111;
12'b000011100000: dataB <= 32'b01101010001101101010010100101011;
12'b000011100001: dataB <= 32'b00000001100111011110000100101011;
12'b000011100010: dataB <= 32'b01000111100001101110111000111000;
12'b000011100011: dataB <= 32'b00000110100101010010011110111011;
12'b000011100100: dataB <= 32'b11010001001011100010000001110100;
12'b000011100101: dataB <= 32'b00000010100101000100101010111010;
12'b000011100110: dataB <= 32'b10100110100101110011000000101110;
12'b000011100111: dataB <= 32'b00000100010001110100010100101100;
12'b000011101000: dataB <= 32'b10011101100011011110011111010100;
12'b000011101001: dataB <= 32'b00001011001100111000100010101111;
12'b000011101010: dataB <= 32'b10100000011000110011100101001010;
12'b000011101011: dataB <= 32'b00001001001010011000110000101011;
12'b000011101100: dataB <= 32'b01010111100010011110011111010000;
12'b000011101101: dataB <= 32'b00000010110111110010100101100111;
12'b000011101110: dataB <= 32'b01001011011101111110110101011100;
12'b000011101111: dataB <= 32'b00000111111110001111110001100101;
12'b000011110000: dataB <= 32'b10011110101101000111001111001011;
12'b000011110001: dataB <= 32'b00000100011101001101101001011011;
12'b000011110010: dataB <= 32'b11100111000101110010100100100010;
12'b000011110011: dataB <= 32'b00001001100010000100101101010101;
12'b000011110100: dataB <= 32'b00110011000101110111011101010101;
12'b000011110101: dataB <= 32'b00001000101000101010010100111111;
12'b000011110110: dataB <= 32'b00100111001001110001110101001001;
12'b000011110111: dataB <= 32'b00001101101101011001010011110101;
12'b000011111000: dataB <= 32'b00010001100010011010100111001101;
12'b000011111001: dataB <= 32'b00001000110001011011001111110011;
12'b000011111010: dataB <= 32'b10011111000001010111011001010101;
12'b000011111011: dataB <= 32'b00000100101001011000001110011011;
12'b000011111100: dataB <= 32'b11010101000101001101101011101110;
12'b000011111101: dataB <= 32'b00001001111010110001010101110011;
12'b000011111110: dataB <= 32'b00010010010010110100010110010101;
12'b000011111111: dataB <= 32'b00001110110110110011000001111001;
12'b000100000000: dataB <= 32'b01011101101111010110101010110100;
12'b000100000001: dataB <= 32'b00001010111110100111011010010110;
12'b000100000010: dataB <= 32'b01101001000111001100111001011000;
12'b000100000011: dataB <= 32'b00000110001000011110000101001111;
12'b000100000100: dataB <= 32'b00000010111001011100000011110100;
12'b000100000101: dataB <= 32'b00000000101010001010011100010011;
12'b000100000110: dataB <= 32'b01010011000011101101111100110000;
12'b000100000111: dataB <= 32'b00000010000110010010010001110011;
12'b000100001000: dataB <= 32'b10011011111000111100010001010011;
12'b000100001001: dataB <= 32'b00001001110011101110111010010111;
12'b000100001010: dataB <= 32'b11100100000100111101011011100111;
12'b000100001011: dataB <= 32'b00000101001110011010100010010000;
12'b000100001100: dataB <= 32'b10100001000010011101100111010111;
12'b000100001101: dataB <= 32'b00000110111110111100111101110101;
12'b000100001110: dataB <= 32'b01110110110000011100000011101100;
12'b000100001111: dataB <= 32'b00000011011001010011010111110011;
12'b000100010000: dataB <= 32'b10101100101011011100111111001101;
12'b000100010001: dataB <= 32'b00000111111110100001100010010011;
12'b000100010010: dataB <= 32'b10011010000110110111010111111101;
12'b000100010011: dataB <= 32'b00000011101100001110010100001100;
12'b000100010100: dataB <= 32'b00011101010010111100000101011000;
12'b000100010101: dataB <= 32'b00000101100010001110010101010110;
12'b000100010110: dataB <= 32'b10010010100111101101010110011010;
12'b000100010111: dataB <= 32'b00001101100110010101000100110011;
12'b000100011000: dataB <= 32'b10110000101101001100110110001110;
12'b000100011001: dataB <= 32'b00000001010100000010111101010110;
12'b000100011010: dataB <= 32'b00000010101101110001010010101100;
12'b000100011011: dataB <= 32'b00001011111101101111011000111011;
12'b000100011100: dataB <= 32'b11100000011011010110101001110110;
12'b000100011101: dataB <= 32'b00000101000001100000000101101010;
12'b000100011110: dataB <= 32'b10011001010111110100010111010010;
12'b000100011111: dataB <= 32'b00000010010110011110101110001100;
12'b000100100000: dataB <= 32'b01010001010011101101111011010110;
12'b000100100001: dataB <= 32'b00000110100101000010111010001011;
12'b000100100010: dataB <= 32'b11001011101011011011100100111100;
12'b000100100011: dataB <= 32'b00000110110110110000110110011011;
12'b000100100100: dataB <= 32'b10111000011101000100001001100001;
12'b000100100101: dataB <= 32'b00001000110111011001101001011101;
12'b000100100110: dataB <= 32'b01001010101011000101011101010000;
12'b000100100111: dataB <= 32'b00001010000101100100000101001011;
12'b000100101000: dataB <= 32'b01101000000101011110110110110110;
12'b000100101001: dataB <= 32'b00001100110000100001010010000001;
12'b000100101010: dataB <= 32'b01000101010000100011100000110001;
12'b000100101011: dataB <= 32'b00000101111110011101101101011011;
12'b000100101100: dataB <= 32'b10100101110001100100010111101101;
12'b000100101101: dataB <= 32'b00000111101000000010101010000111;
12'b000100101110: dataB <= 32'b00101010101100010101001010100001;
12'b000100101111: dataB <= 32'b00001011001100100000110111100010;
12'b000100110000: dataB <= 32'b11010001000101011011111001100110;
12'b000100110001: dataB <= 32'b00001010110110101111000100010101;
12'b000100110010: dataB <= 32'b01011010111110001110001001110010;
12'b000100110011: dataB <= 32'b00001111010001001011101000111110;
12'b000100110100: dataB <= 32'b10110001001010000011100010010101;
12'b000100110101: dataB <= 32'b00000110111000100001010010000111;
12'b000100110110: dataB <= 32'b11100110001001100010010100001101;
12'b000100110111: dataB <= 32'b00000001001010011000001000101011;
12'b000100111000: dataB <= 32'b00001011101001111111001001011000;
12'b000100111001: dataB <= 32'b00000101100110001110100010111011;
12'b000100111010: dataB <= 32'b10010011010011010001010010010110;
12'b000100111011: dataB <= 32'b00000001101000000010110110110010;
12'b000100111100: dataB <= 32'b00100100100101101011000000110001;
12'b000100111101: dataB <= 32'b00000100110010110000001100110101;
12'b000100111110: dataB <= 32'b00100001100011101101111111010001;
12'b000100111111: dataB <= 32'b00001010101011110100010110111111;
12'b000101000000: dataB <= 32'b01011100011000110100000101001011;
12'b000101000001: dataB <= 32'b00001000101001011000110000101100;
12'b000101000010: dataB <= 32'b01011001100010101110001111001101;
12'b000101000011: dataB <= 32'b00000011011001101110100001111111;
12'b000101000100: dataB <= 32'b10001111100110001110110110011101;
12'b000101000101: dataB <= 32'b00001001011110010101110101101101;
12'b000101000110: dataB <= 32'b11011110101101011111101110101000;
12'b000101000111: dataB <= 32'b00000101111110010011110001011011;
12'b000101001000: dataB <= 32'b00100111000101100010100011100011;
12'b000101001001: dataB <= 32'b00001000000010000010111001100110;
12'b000101001010: dataB <= 32'b01110010111110000111011101010011;
12'b000101001011: dataB <= 32'b00001000001000100110010001010111;
12'b000101001100: dataB <= 32'b01101001000101101001110100101011;
12'b000101001101: dataB <= 32'b00001101001011011011010011110100;
12'b000101001110: dataB <= 32'b01010101101010010010010111001101;
12'b000101001111: dataB <= 32'b00001001010000011101010011101010;
12'b000101010000: dataB <= 32'b10011111000001101111101001110100;
12'b000101010001: dataB <= 32'b00000100001010010100010010011011;
12'b000101010010: dataB <= 32'b11010101001101010110001011001101;
12'b000101010011: dataB <= 32'b00001010111001110011001101110011;
12'b000101010100: dataB <= 32'b01001110010110110011110110110110;
12'b000101010101: dataB <= 32'b00001111010011110010111001101001;
12'b000101010110: dataB <= 32'b00100001101111100110001011010011;
12'b000101010111: dataB <= 32'b00001011111100101001010110100110;
12'b000101011000: dataB <= 32'b10101001000011010100011010010111;
12'b000101011001: dataB <= 32'b00000101101001011010001001100111;
12'b000101011010: dataB <= 32'b11000011000101011100010100010110;
12'b000101011011: dataB <= 32'b00000000101101001000101000010011;
12'b000101011100: dataB <= 32'b10010011000111110101001100101111;
12'b000101011101: dataB <= 32'b00000001001000001110011001101011;
12'b000101011110: dataB <= 32'b01100001111000111100110001110110;
12'b000101011111: dataB <= 32'b00001010010010101110110110101111;
12'b000101100000: dataB <= 32'b11011110000101000101111010100110;
12'b000101100001: dataB <= 32'b00000101001111011000100110000000;
12'b000101100010: dataB <= 32'b10100001000010100101011000010111;
12'b000101100011: dataB <= 32'b00001000011110111010110101111101;
12'b000101100100: dataB <= 32'b10110100101000100100110011001110;
12'b000101100101: dataB <= 32'b00000100011010010101011011110010;
12'b000101100110: dataB <= 32'b10101010100111100100001110101010;
12'b000101100111: dataB <= 32'b00001001011110100101100010010011;
12'b000101101000: dataB <= 32'b01010110000111000111001001011101;
12'b000101101001: dataB <= 32'b00000011101110001010011100010101;
12'b000101101010: dataB <= 32'b01011111010010111011100101111001;
12'b000101101011: dataB <= 32'b00000100100011001010011101011110;
12'b000101101100: dataB <= 32'b00010000101111110100100111011011;
12'b000101101101: dataB <= 32'b00001100100100010111001000110100;
12'b000101101110: dataB <= 32'b11101110101001010101000110001111;
12'b000101101111: dataB <= 32'b00000001110110000011001001100110;
12'b000101110000: dataB <= 32'b10000010111001100001010010101110;
12'b000101110001: dataB <= 32'b00001100111011110001010000111011;
12'b000101110010: dataB <= 32'b00011100011011100101111010010101;
12'b000101110011: dataB <= 32'b00000100000011011010000101100011;
12'b000101110100: dataB <= 32'b01011011010111110011100111010010;
12'b000101110101: dataB <= 32'b00000011011000011100101110010100;
12'b000101110110: dataB <= 32'b01010011011011110101001011110100;
12'b000101110111: dataB <= 32'b00000101100101000011000110001011;
12'b000101111000: dataB <= 32'b10010001110011010011000101111101;
12'b000101111001: dataB <= 32'b00000111110111101110101110011011;
12'b000101111010: dataB <= 32'b11110100010101001100101000000001;
12'b000101111011: dataB <= 32'b00001001010111011101101001100101;
12'b000101111100: dataB <= 32'b11001000110011000100111101001110;
12'b000101111101: dataB <= 32'b00001001000101011110000101000011;
12'b000101111110: dataB <= 32'b01100010000101101111000111110111;
12'b000101111111: dataB <= 32'b00001100101110100011010001110001;
12'b000110000000: dataB <= 32'b10000111011000100100010000110100;
12'b000110000001: dataB <= 32'b00000111011110100011101101010011;
12'b000110000010: dataB <= 32'b10101001101101100100100111101101;
12'b000110000011: dataB <= 32'b00000110101001000010110110011111;
12'b000110000100: dataB <= 32'b01101000101000011101101001000001;
12'b000110000101: dataB <= 32'b00001010101011100000110111010001;
12'b000110000110: dataB <= 32'b01010001001001011100001000100101;
12'b000110000111: dataB <= 32'b00001011010101101110111100100110;
12'b000110001000: dataB <= 32'b11011011000010011110001001110001;
12'b000110001001: dataB <= 32'b00001111001110010001110001001110;
12'b000110001010: dataB <= 32'b10110001000001111011100010111000;
12'b000110001011: dataB <= 32'b00000111111000100011010010011111;
12'b000110001100: dataB <= 32'b01100000001001011010100100001110;
12'b000110001101: dataB <= 32'b00000000101101010010001100101100;
12'b000110001110: dataB <= 32'b11010001110010001110111010010111;
12'b000110001111: dataB <= 32'b00000101000111001100101010110010;
12'b000110010000: dataB <= 32'b01010101010111000000110011011000;
12'b000110010001: dataB <= 32'b00000000101010000011000010101010;
12'b000110010010: dataB <= 32'b01100000100001100011010000110100;
12'b000110010011: dataB <= 32'b00000101010100101100001000111101;
12'b000110010100: dataB <= 32'b10100101100011110101001111001110;
12'b000110010101: dataB <= 32'b00001010001010110000001111010110;
12'b000110010110: dataB <= 32'b11011000011100110100100100101101;
12'b000110010111: dataB <= 32'b00001000001001010110110100101100;
12'b000110011000: dataB <= 32'b01011101100110111101111111001010;
12'b000110011001: dataB <= 32'b00000100011010101100011010010111;
12'b000110011010: dataB <= 32'b10010011101110011110100111111101;
12'b000110011011: dataB <= 32'b00001010111110011011111001110101;
12'b000110011100: dataB <= 32'b00011100101101101111101101100110;
12'b000110011101: dataB <= 32'b00000111011110010111110101011100;
12'b000110011110: dataB <= 32'b00100111000001011010110010100101;
12'b000110011111: dataB <= 32'b00000110100010000011000101110110;
12'b000110100000: dataB <= 32'b10110010110110011111011101110001;
12'b000110100001: dataB <= 32'b00000111001000100000001101101111;
12'b000110100010: dataB <= 32'b10101001000001011010000100001100;
12'b000110100011: dataB <= 32'b00001100101001011101010111110011;
12'b000110100100: dataB <= 32'b11011001101110001010010110101110;
12'b000110100101: dataB <= 32'b00001001010000011111010011100001;
12'b000110100110: dataB <= 32'b01011111000010000111101010010011;
12'b000110100111: dataB <= 32'b00000011101011001110010110011011;
12'b000110101000: dataB <= 32'b00010111010001100110001010101011;
12'b000110101001: dataB <= 32'b00001011111000110101000101110100;
12'b000110101010: dataB <= 32'b01001010011110110011100111010110;
12'b000110101011: dataB <= 32'b00001111010000110000110001011001;
12'b000110101100: dataB <= 32'b11100101101111101101101011110010;
12'b000110101101: dataB <= 32'b00001101011010101011010010110101;
12'b000110101110: dataB <= 32'b10101001000011010011111010110110;
12'b000110101111: dataB <= 32'b00000100101010010100001001111111;
12'b000110110000: dataB <= 32'b01000011010001100100100100110111;
12'b000110110001: dataB <= 32'b00000000110000000110110000010100;
12'b000110110010: dataB <= 32'b10010101001011110100011100101101;
12'b000110110011: dataB <= 32'b00000000101011001010100001101011;
12'b000110110100: dataB <= 32'b00100111111001000101010010011000;
12'b000110110101: dataB <= 32'b00001010010001101100101111000111;
12'b000110110110: dataB <= 32'b11011000000101010110001001100101;
12'b000110110111: dataB <= 32'b00000101010000010110101001101000;
12'b000110111000: dataB <= 32'b10100001000010101101001000110111;
12'b000110111001: dataB <= 32'b00001001111110111010101010001101;
12'b000110111010: dataB <= 32'b00110000100000101101010011010000;
12'b000110111011: dataB <= 32'b00000101011011011001011111100010;
12'b000110111100: dataB <= 32'b01101000100011100011101110000111;
12'b000110111101: dataB <= 32'b00001010011110100111011110010011;
12'b000110111110: dataB <= 32'b00010000001111010110101010011100;
12'b000110111111: dataB <= 32'b00000011101111001000100100011110;
12'b000111000000: dataB <= 32'b10011111010010111011010110111010;
12'b000111000001: dataB <= 32'b00000011000101001000100101101110;
12'b000111000010: dataB <= 32'b01001110110011110100001000011011;
12'b000111000011: dataB <= 32'b00001011100010010111001100110100;
12'b000111000100: dataB <= 32'b00101100100101011101010110010000;
12'b000111000101: dataB <= 32'b00000010111001000101010101111111;
12'b000111000110: dataB <= 32'b11000011000101010001100010110001;
12'b000111000111: dataB <= 32'b00001101111001110011001000111011;
12'b000111001000: dataB <= 32'b00011000011111110101011010110100;
12'b000111001001: dataB <= 32'b00000010100101010100001001100011;
12'b000111001010: dataB <= 32'b01011101011011110010110111110011;
12'b000111001011: dataB <= 32'b00000100011010011010101110010100;
12'b000111001100: dataB <= 32'b00010101011111110100011100010011;
12'b000111001101: dataB <= 32'b00000100100110000011010010000011;
12'b000111001110: dataB <= 32'b10010101111011010010100111011101;
12'b000111001111: dataB <= 32'b00001000010111101100101010011011;
12'b000111010000: dataB <= 32'b11101110001101001100110110100001;
12'b000111010001: dataB <= 32'b00001010010110100011101001101101;
12'b000111010010: dataB <= 32'b00000110111111001100011100101100;
12'b000111010011: dataB <= 32'b00001000000100011000000101000100;
12'b000111010100: dataB <= 32'b10011100000110000111001000010111;
12'b000111010101: dataB <= 32'b00001100001100100101001101100001;
12'b000111010110: dataB <= 32'b11001011100100101100110001010110;
12'b000111010111: dataB <= 32'b00001000111110100111101001010011;
12'b000111011000: dataB <= 32'b01101101101001101100110111001110;
12'b000111011001: dataB <= 32'b00000110001001000011000010110111;
12'b000111011010: dataB <= 32'b11100110100100101110010111100001;
12'b000111011011: dataB <= 32'b00001010001010100000110111000000;
12'b000111011100: dataB <= 32'b11010011010001011100010111100101;
12'b000111011101: dataB <= 32'b00001011110011101110111000110110;
12'b000111011110: dataB <= 32'b00011011000010101101111001110001;
12'b000111011111: dataB <= 32'b00001111001011010101111001011111;
12'b000111100000: dataB <= 32'b01110000111001111011100011111010;
12'b000111100001: dataB <= 32'b00001000111000100101001110110111;
12'b000111100010: dataB <= 32'b11011100001001010010110011110000;
12'b000111100011: dataB <= 32'b00000000101111001110010000110100;
12'b000111100100: dataB <= 32'b01010101111010100110111010110110;
12'b000111100101: dataB <= 32'b00000100001000001010110010101010;
12'b000111100110: dataB <= 32'b00010111011010110000100100011010;
12'b000111100111: dataB <= 32'b00000000101101000011001110100010;
12'b000111101000: dataB <= 32'b11011110100001100011100001010110;
12'b000111101001: dataB <= 32'b00000101010101100110000101000101;
12'b000111101010: dataB <= 32'b00100111011111110100011111001011;
12'b000111101011: dataB <= 32'b00001001101001101100001011100110;
12'b000111101100: dataB <= 32'b01010110011100110101000100001110;
12'b000111101101: dataB <= 32'b00000111001001010110111000110101;
12'b000111101110: dataB <= 32'b00100001100111000101011110001000;
12'b000111101111: dataB <= 32'b00000101011011101000010110100111;
12'b000111110000: dataB <= 32'b10010111110010101110101000111101;
12'b000111110001: dataB <= 32'b00001011111100100001111001111101;
12'b000111110010: dataB <= 32'b01011010110010000111101100100100;
12'b000111110011: dataB <= 32'b00001000111110011101110101011100;
12'b000111110100: dataB <= 32'b00100110111101011011000001101000;
12'b000111110101: dataB <= 32'b00000101100011000101010001111110;
12'b000111110110: dataB <= 32'b10110010101110101111001101101111;
12'b000111110111: dataB <= 32'b00000110101000011100001101111111;
12'b000111111000: dataB <= 32'b11101001000001010010010100001101;
12'b000111111001: dataB <= 32'b00001011100111011111010111110010;
12'b000111111010: dataB <= 32'b01011101101110000010010110101110;
12'b000111111011: dataB <= 32'b00001001010000011111010011010001;
12'b000111111100: dataB <= 32'b00011111000010011111101010110010;
12'b000111111101: dataB <= 32'b00000011101101001010011110010011;
12'b000111111110: dataB <= 32'b00011001010001110110011010101010;
12'b000111111111: dataB <= 32'b00001100010110110100111101110100;
12'b001000000000: dataB <= 32'b10001000100110101011010111110110;
12'b001000000001: dataB <= 32'b00001111001101110000101101001001;
12'b001000000010: dataB <= 32'b10101001101011110100111011110000;
12'b001000000011: dataB <= 32'b00001110011000101101001110111101;
12'b001000000100: dataB <= 32'b10101000111111010011011011010101;
12'b001000000101: dataB <= 32'b00000100001011010000010010010111;
12'b001000000110: dataB <= 32'b00000101011101100100110101111000;
12'b001000000111: dataB <= 32'b00000000110011000100111100011101;
12'b001000001000: dataB <= 32'b11010101001111110011101100001011;
12'b001000001001: dataB <= 32'b00000000101110001000101001101011;
12'b001000001010: dataB <= 32'b10101011110101001101100011011010;
12'b001000001011: dataB <= 32'b00001010110000101010101011010110;
12'b001000001100: dataB <= 32'b00010010001001100110011000100100;
12'b001000001101: dataB <= 32'b00000101010001010100101101011001;
12'b001000001110: dataB <= 32'b01100001000010110100101001110111;
12'b001000001111: dataB <= 32'b00001010111101110110100010010101;
12'b001000010000: dataB <= 32'b01101110011000110101110011010010;
12'b001000010001: dataB <= 32'b00000110111100011011011111011001;
12'b001000010010: dataB <= 32'b01100100011111011011001101000101;
12'b001000010011: dataB <= 32'b00001011111100101011011010001011;
12'b001000010100: dataB <= 32'b10001100010011100101111011011011;
12'b001000010101: dataB <= 32'b00000011110001000110110000101110;
12'b001000010110: dataB <= 32'b10100001010010110010110111111010;
12'b001000010111: dataB <= 32'b00000010100111000110110001111110;
12'b001000011000: dataB <= 32'b11001110111011110011011001011011;
12'b001000011001: dataB <= 32'b00001010000001011001010000111100;
12'b001000011010: dataB <= 32'b11101000011101101101100110010001;
12'b001000011011: dataB <= 32'b00000011111010000111100010001110;
12'b001000011100: dataB <= 32'b01000011010001001001110010110011;
12'b001000011101: dataB <= 32'b00001110110111110101000000111100;
12'b001000011110: dataB <= 32'b01010110100011110100101011010010;
12'b001000011111: dataB <= 32'b00000001100111001110001101011011;
12'b001000100000: dataB <= 32'b00100001011011101010001000010011;
12'b001000100001: dataB <= 32'b00000101011011011010101110010100;
12'b001000100010: dataB <= 32'b00011001100011110011101100010001;
12'b001000100011: dataB <= 32'b00000011101000000101011101111011;
12'b001000100100: dataB <= 32'b01011011111011000010001000111101;
12'b001000100101: dataB <= 32'b00001001010110101010100110010011;
12'b001000100110: dataB <= 32'b00101010000101010101000101100001;
12'b001000100111: dataB <= 32'b00001010110101100111101001111110;
12'b001000101000: dataB <= 32'b10001001000111001011111100101010;
12'b001000101001: dataB <= 32'b00000111000100010010001001001100;
12'b001000101010: dataB <= 32'b10010110000110010111001001010110;
12'b001000101011: dataB <= 32'b00001011101011100111001101010001;
12'b001000101100: dataB <= 32'b00001111101000110101010010011001;
12'b001000101101: dataB <= 32'b00001010011110101011100101010100;
12'b001000101110: dataB <= 32'b11110001100001101100110111001110;
12'b001000101111: dataB <= 32'b00000101101010000011001111001110;
12'b001000110000: dataB <= 32'b10100100100100111110100110000001;
12'b001000110001: dataB <= 32'b00001001001001011110110110110000;
12'b001000110010: dataB <= 32'b01010101010101100100010110100101;
12'b001000110011: dataB <= 32'b00001011110010101110110001000111;
12'b001000110100: dataB <= 32'b01011011000110110101101010010000;
12'b001000110101: dataB <= 32'b00001110101000011011111001110111;
12'b001000110110: dataB <= 32'b11110000110101111011100100111011;
12'b001000110111: dataB <= 32'b00001001011000100111001111001110;
12'b001000111000: dataB <= 32'b01010110001101001011010100010001;
12'b001000111001: dataB <= 32'b00000000110010001010011000110101;
12'b001000111010: dataB <= 32'b00011011111010110110101011010101;
12'b001000111011: dataB <= 32'b00000011101010001000111010100010;
12'b001000111100: dataB <= 32'b11011001011110011000010101011011;
12'b001000111101: dataB <= 32'b00000000110000000101010110010001;
12'b001000111110: dataB <= 32'b00011010100101100011100010011001;
12'b001000111111: dataB <= 32'b00000110010110100000000101010110;
12'b001001000000: dataB <= 32'b10101011011011110011101110101000;
12'b001001000001: dataB <= 32'b00001001001001100110000111101101;
12'b001001000010: dataB <= 32'b10010010100000111101010100001111;
12'b001001000011: dataB <= 32'b00000110101010010100111100111101;
12'b001001000100: dataB <= 32'b11100101100111001100111101100101;
12'b001001000101: dataB <= 32'b00000110111100100100010110110110;
12'b001001000110: dataB <= 32'b10011101110110111110001010011100;
12'b001001000111: dataB <= 32'b00001101011011100101111010001101;
12'b001001001000: dataB <= 32'b01011000110010011111101011100010;
12'b001001001001: dataB <= 32'b00001010011110100011110101100100;
12'b001001001010: dataB <= 32'b00100110111001010011010000101010;
12'b001001001011: dataB <= 32'b00000100100100000111011010001110;
12'b001001001100: dataB <= 32'b10110000101011000110101101101101;
12'b001001001101: dataB <= 32'b00000101101001011000010010010111;
12'b001001001110: dataB <= 32'b00101000111101001010100011101111;
12'b001001001111: dataB <= 32'b00001011000110100001010111101010;
12'b001001010000: dataB <= 32'b11100001101101110010010110101111;
12'b001001010001: dataB <= 32'b00001001001111100001010010111000;
12'b001001010010: dataB <= 32'b00011111000010101111011010110001;
12'b001001010011: dataB <= 32'b00000011001111001000100110010011;
12'b001001010100: dataB <= 32'b00011011010110000110011001101001;
12'b001001010101: dataB <= 32'b00001100110101110100110101110100;
12'b001001010110: dataB <= 32'b00000110110010101011001000110110;
12'b001001010111: dataB <= 32'b00001111001011101110100100111010;
12'b001001011000: dataB <= 32'b00101101100111110100001011101111;
12'b001001011001: dataB <= 32'b00001110110110101101001011000101;
12'b001001011010: dataB <= 32'b10101000111011001010111011110011;
12'b001001011011: dataB <= 32'b00000100001101001010010110100111;
12'b001001011100: dataB <= 32'b10001001100101101100110110111001;
12'b001001011101: dataB <= 32'b00000001010110000101000100100101;
12'b001001011110: dataB <= 32'b11010111010011110010111011101001;
12'b001001011111: dataB <= 32'b00000000110001000110110001101011;
12'b001001100000: dataB <= 32'b00110001110001011101110100011100;
12'b001001100001: dataB <= 32'b00001010101111101000100111100110;
12'b001001100010: dataB <= 32'b01001110001101110110010111100100;
12'b001001100011: dataB <= 32'b00000101010010010010110001001001;
12'b001001100100: dataB <= 32'b01100001000010110100011010010110;
12'b001001100101: dataB <= 32'b00001100011100110100010110011101;
12'b001001100110: dataB <= 32'b11101010010101000110010011110100;
12'b001001100111: dataB <= 32'b00000111111101011111011111000000;
12'b001001101000: dataB <= 32'b01100000011111010010101100000011;
12'b001001101001: dataB <= 32'b00001100111011101101010110001011;
12'b001001101010: dataB <= 32'b00001000011011110101011100111001;
12'b001001101011: dataB <= 32'b00000011110011000110111000111111;
12'b001001101100: dataB <= 32'b10100011010010101010101001011010;
12'b001001101101: dataB <= 32'b00000001101001000110111010010110;
12'b001001101110: dataB <= 32'b01001101000011101010101010011010;
12'b001001101111: dataB <= 32'b00001000100001011011010001000101;
12'b001001110000: dataB <= 32'b11100100011101110101100110010001;
12'b001001110001: dataB <= 32'b00000100111100001011101010011110;
12'b001001110010: dataB <= 32'b11000101011100111010010011010101;
12'b001001110011: dataB <= 32'b00001111010100110100111000111100;
12'b001001110100: dataB <= 32'b10010010100111110011111011010001;
12'b001001110101: dataB <= 32'b00000001001001001010010101011011;
12'b001001110110: dataB <= 32'b00100011011011011001101000010011;
12'b001001110111: dataB <= 32'b00000110011100011000110010010100;
12'b001001111000: dataB <= 32'b00011101100011110010111100101111;
12'b001001111001: dataB <= 32'b00000011001010001001100101111011;
12'b001001111010: dataB <= 32'b01100001111010110001101001111101;
12'b001001111011: dataB <= 32'b00001001110110100110100010010011;
12'b001001111100: dataB <= 32'b00100100000101011101010100000011;
12'b001001111101: dataB <= 32'b00001011010100101011100110001110;
12'b001001111110: dataB <= 32'b11001001001111001011011011101000;
12'b001001111111: dataB <= 32'b00000110000101001110010001001100;
12'b001010000000: dataB <= 32'b00010000001010100110111001110110;
12'b001010000001: dataB <= 32'b00001011001001100111001001000010;
12'b001010000010: dataB <= 32'b01010011110000111101110011011011;
12'b001010000011: dataB <= 32'b00001011111101101111100001010100;
12'b001010000100: dataB <= 32'b10110101011101110100110111001110;
12'b001010000101: dataB <= 32'b00000101001011000101011011011110;
12'b001010000110: dataB <= 32'b01100000100101001111000100100010;
12'b001010000111: dataB <= 32'b00001000101001011110110110011000;
12'b001010001000: dataB <= 32'b10010111011001100100100101100110;
12'b001010001001: dataB <= 32'b00001011110000101100101101011111;
12'b001010001010: dataB <= 32'b01011011000110111101001010001111;
12'b001010001011: dataB <= 32'b00001101100110100001111010000111;
12'b001010001100: dataB <= 32'b10101110101101111011100101111100;
12'b001010001101: dataB <= 32'b00001010010111100111001011011110;
12'b001010001110: dataB <= 32'b11010010010001001011100100010011;
12'b001010001111: dataB <= 32'b00000001010101000110100001000101;
12'b001010010000: dataB <= 32'b00100001111011000110001011110011;
12'b001010010001: dataB <= 32'b00000011001100001001000010010010;
12'b001010010010: dataB <= 32'b11011101011110000000010110011100;
12'b001010010011: dataB <= 32'b00000000110011000111100010000001;
12'b001010010100: dataB <= 32'b01011000100101100011110011011011;
12'b001010010101: dataB <= 32'b00000110110110011010000101100110;
12'b001010010110: dataB <= 32'b11101101010111110010111101100110;
12'b001010010111: dataB <= 32'b00001000001001100000000111110100;
12'b001010011000: dataB <= 32'b00010000101001001101110100010001;
12'b001010011001: dataB <= 32'b00000110001010010101000001001110;
12'b001010011010: dataB <= 32'b01101001100011001100011100000011;
12'b001010011011: dataB <= 32'b00000111111101100000010011001110;
12'b001010011100: dataB <= 32'b10100001110111001101101011011011;
12'b001010011101: dataB <= 32'b00001110011000101011110110010101;
12'b001010011110: dataB <= 32'b10011000110110110111011010000001;
12'b001010011111: dataB <= 32'b00001011111101100111110101100100;
12'b001010100000: dataB <= 32'b00100110111001010011100000101101;
12'b001010100001: dataB <= 32'b00000011000110001011100010011110;
12'b001010100010: dataB <= 32'b01101100100011010110011101001011;
12'b001010100011: dataB <= 32'b00000101001010010100010110101111;
12'b001010100100: dataB <= 32'b10101000111001000011000011110001;
12'b001010100101: dataB <= 32'b00001010000101100011010111011001;
12'b001010100110: dataB <= 32'b01100101101101101010010110101111;
12'b001010100111: dataB <= 32'b00001001001111100011010010101000;
12'b001010101000: dataB <= 32'b00011111000011000111001010110000;
12'b001010101001: dataB <= 32'b00000011010001000110101110001011;
12'b001010101010: dataB <= 32'b00011101010110010110011001001001;
12'b001010101011: dataB <= 32'b00001101010011110010101101110100;
12'b001010101100: dataB <= 32'b10000110111010100010111001010110;
12'b001010101101: dataB <= 32'b00001110001000101010100000110010;
12'b001010101110: dataB <= 32'b10110001011111110011011011101101;
12'b001010101111: dataB <= 32'b00001111010011101101000011001100;
12'b001010110000: dataB <= 32'b11011100101101011001101001101000;
12'b001010110001: dataB <= 32'b00000110110111001011101011110010;
12'b001010110010: dataB <= 32'b11110011101110011100101100110010;
12'b001010110011: dataB <= 32'b00001011011101100011110110110110;
12'b001010110100: dataB <= 32'b10101001010001011000010100101000;
12'b001010110101: dataB <= 32'b00001000111110011001110001111100;
12'b001010110110: dataB <= 32'b11111000011110111101001110010111;
12'b001010110111: dataB <= 32'b00000111101010010010101111000000;
12'b001010111000: dataB <= 32'b10000111100011001100010010010000;
12'b001010111001: dataB <= 32'b00001001010101011001011000101101;
12'b001010111010: dataB <= 32'b00100000111110001010011011001011;
12'b001010111011: dataB <= 32'b00001110000111001010010110101011;
12'b001010111100: dataB <= 32'b11001010101011001101111010011000;
12'b001010111101: dataB <= 32'b00001110110000101111000000011001;
12'b001010111110: dataB <= 32'b10001110111101010001010001100111;
12'b001010111111: dataB <= 32'b00001101100110101010100101101011;
12'b001011000000: dataB <= 32'b00001101101110101000011100100110;
12'b001011000001: dataB <= 32'b00001001111000011101110011100110;
12'b001011000010: dataB <= 32'b01101000111001010010101101001101;
12'b001011000011: dataB <= 32'b00000100111100011101110011010011;
12'b001011000100: dataB <= 32'b11100001100101010000101101001011;
12'b001011000101: dataB <= 32'b00000000101110101001001010101101;
12'b001011000110: dataB <= 32'b00001110110110110100011000110011;
12'b001011000111: dataB <= 32'b00001110010110110101101011011011;
12'b001011001000: dataB <= 32'b00101111110101001110001010111001;
12'b001011001001: dataB <= 32'b00001010000001011100010110011110;
12'b001011001010: dataB <= 32'b00010011011001111000011000101001;
12'b001011001011: dataB <= 32'b00000100111101001011101001110101;
12'b001011001100: dataB <= 32'b01101100111000110001001001101111;
12'b001011001101: dataB <= 32'b00001110010011011001001110000011;
12'b001011001110: dataB <= 32'b00110001000101011000010111100110;
12'b001011001111: dataB <= 32'b00000101011001110011101101100100;
12'b001011010000: dataB <= 32'b01111100111100110010011110101100;
12'b001011010001: dataB <= 32'b00001011001100010000110001101011;
12'b001011010010: dataB <= 32'b10000010110110101101000001110111;
12'b001011010011: dataB <= 32'b00001010001001110010101011000011;
12'b001011010100: dataB <= 32'b10100111101101101001100100001000;
12'b001011010101: dataB <= 32'b00000010110011001001100010011101;
12'b001011010110: dataB <= 32'b11000101011111011010111011001100;
12'b001011010111: dataB <= 32'b00000100101001100100110001000101;
12'b001011011000: dataB <= 32'b01111001011010111110001101111001;
12'b001011011001: dataB <= 32'b00001110101000110000100010001101;
12'b001011011010: dataB <= 32'b00101110010110011100010111010001;
12'b001011011011: dataB <= 32'b00000101110101101101110111010001;
12'b001011011100: dataB <= 32'b00010010111111100101100001010110;
12'b001011011101: dataB <= 32'b00000100101110011011000000001011;
12'b001011011110: dataB <= 32'b00101101010010010100110011010100;
12'b001011011111: dataB <= 32'b00001000001000010110100111110101;
12'b001011100000: dataB <= 32'b11100011001010100010000111101011;
12'b001011100001: dataB <= 32'b00000011000100111100111111101011;
12'b001011100010: dataB <= 32'b00010110100001110100001110010100;
12'b001011100011: dataB <= 32'b00001011101011100100110011010001;
12'b001011100100: dataB <= 32'b11001001011001110101101001110111;
12'b001011100101: dataB <= 32'b00001010111101010001110010111101;
12'b001011100110: dataB <= 32'b01111100111111000001111001101000;
12'b001011100111: dataB <= 32'b00000110011001100001101101000011;
12'b001011101000: dataB <= 32'b11101111000100001011111110010011;
12'b001011101001: dataB <= 32'b00001001111110110001110000111011;
12'b001011101010: dataB <= 32'b11010011001101111100111101111001;
12'b001011101011: dataB <= 32'b00001011010010000011001011001100;
12'b001011101100: dataB <= 32'b01101010100101011000010011000100;
12'b001011101101: dataB <= 32'b00000100101111000010111110011000;
12'b001011101110: dataB <= 32'b10010101011110111101101000110111;
12'b001011101111: dataB <= 32'b00000101010011100001010111000101;
12'b001011110000: dataB <= 32'b10110000101110001001100001100111;
12'b001011110001: dataB <= 32'b00001110110000001000111111001001;
12'b001011110010: dataB <= 32'b01111010111110110001101101101001;
12'b001011110011: dataB <= 32'b00001100000011111010101010110011;
12'b001011110100: dataB <= 32'b11011011001111101010010000101011;
12'b001011110101: dataB <= 32'b00001110101000111010110010010100;
12'b001011110110: dataB <= 32'b00011100110001110101010110111110;
12'b001011110111: dataB <= 32'b00000011011001110001101011000011;
12'b001011111000: dataB <= 32'b10010000100111001001010101100101;
12'b001011111001: dataB <= 32'b00000101010101001011010111101010;
12'b001011111010: dataB <= 32'b00011100101101100101111000111000;
12'b001011111011: dataB <= 32'b00000010101011101010111000110001;
12'b001011111100: dataB <= 32'b10110110110101001100100111110010;
12'b001011111101: dataB <= 32'b00000111101101101000111000001010;
12'b001011111110: dataB <= 32'b10100001000011100001111000001010;
12'b001011111111: dataB <= 32'b00001000111001010111110001100011;
12'b001100000000: dataB <= 32'b01101011000111001011010100101101;
12'b001100000001: dataB <= 32'b00001001100101010110011010000100;
12'b001100000010: dataB <= 32'b01011101110001011010111011001101;
12'b001100000011: dataB <= 32'b00000100000011010000101001010110;
12'b001100000100: dataB <= 32'b10101110011101101000010110101000;
12'b001100000101: dataB <= 32'b00001001100001100000100110010001;
12'b001100000110: dataB <= 32'b01011110101101101001011010101001;
12'b001100000111: dataB <= 32'b00000101110111001001011111110011;
12'b001100001000: dataB <= 32'b00101111110110011100111100010100;
12'b001100001001: dataB <= 32'b00001001111110011111110110100111;
12'b001100001010: dataB <= 32'b10100111010101110000010101100111;
12'b001100001011: dataB <= 32'b00000111011110010101101101111100;
12'b001100001100: dataB <= 32'b01111010101010110101101101011001;
12'b001100001101: dataB <= 32'b00001000001010010100101011010001;
12'b001100001110: dataB <= 32'b00000101011011001100110010001110;
12'b001100001111: dataB <= 32'b00001000110101010111010100100101;
12'b001100010000: dataB <= 32'b01100000111110010010011011101100;
12'b001100010001: dataB <= 32'b00001110101010010000010010101011;
12'b001100010010: dataB <= 32'b00001100100010111110011001011001;
12'b001100010011: dataB <= 32'b00001110010010101111001000101001;
12'b001100010100: dataB <= 32'b10001110110101100001000010100101;
12'b001100010101: dataB <= 32'b00001110001000101100101001101011;
12'b001100010110: dataB <= 32'b10001001100110111000111101101001;
12'b001100010111: dataB <= 32'b00001000111000011001110011010110;
12'b001100011000: dataB <= 32'b00101000111101011010011101010000;
12'b001100011001: dataB <= 32'b00000011111010011001110011010100;
12'b001100011010: dataB <= 32'b00011101100001101000011101101101;
12'b001100011011: dataB <= 32'b00000000101011101001001110011110;
12'b001100011100: dataB <= 32'b10001110101110110100101000110011;
12'b001100011101: dataB <= 32'b00001101011000110001110011011011;
12'b001100011110: dataB <= 32'b00101001111000111101101001111010;
12'b001100011111: dataB <= 32'b00001011100010100000010110001110;
12'b001100100000: dataB <= 32'b00010001010010010000011001001001;
12'b001100100001: dataB <= 32'b00000011111100000111100001101101;
12'b001100100010: dataB <= 32'b01101100111101000000101001101111;
12'b001100100011: dataB <= 32'b00001101110101010111001010000011;
12'b001100100100: dataB <= 32'b00110001001101110000011000100111;
12'b001100100101: dataB <= 32'b00000100011000101111110101100100;
12'b001100100110: dataB <= 32'b01111101001001000001111110101110;
12'b001100100111: dataB <= 32'b00001011001101010010101001101011;
12'b001100101000: dataB <= 32'b00000010101010100101010000110100;
12'b001100101001: dataB <= 32'b00001010101010110100110011000100;
12'b001100101010: dataB <= 32'b10100011101101111001100101000110;
12'b001100101011: dataB <= 32'b00000010010001000101011010010101;
12'b001100101100: dataB <= 32'b01000011010011100011011011001101;
12'b001100101101: dataB <= 32'b00000101101000100110110000110101;
12'b001100101110: dataB <= 32'b01110101100010101110011100111011;
12'b001100101111: dataB <= 32'b00001111001011110010101010000101;
12'b001100110000: dataB <= 32'b10110000011110011100100111010001;
12'b001100110001: dataB <= 32'b00000101010100100111111011011001;
12'b001100110010: dataB <= 32'b01010010110111010110000000110011;
12'b001100110011: dataB <= 32'b00000100101101011011000000010010;
12'b001100110100: dataB <= 32'b11101011010110001100110010110010;
12'b001100110101: dataB <= 32'b00001001001000011000100011101101;
12'b001100110110: dataB <= 32'b01100011001010110010011000001011;
12'b001100110111: dataB <= 32'b00000100000010111101001011101100;
12'b001100111000: dataB <= 32'b10011010011101110100001101110110;
12'b001100111001: dataB <= 32'b00001100001101100110110011011001;
12'b001100111010: dataB <= 32'b01000111010001101101101000110111;
12'b001100111011: dataB <= 32'b00001001011110001101101010101110;
12'b001100111100: dataB <= 32'b11111101001011010010011010101001;
12'b001100111101: dataB <= 32'b00000101011000011101101101000010;
12'b001100111110: dataB <= 32'b01101111001100001011001101110101;
12'b001100111111: dataB <= 32'b00001000011110101011110100111011;
12'b001101000000: dataB <= 32'b01010011001001110100111100111011;
12'b001101000001: dataB <= 32'b00001011010011000010111111000101;
12'b001101000010: dataB <= 32'b10101100101001110000010100000010;
12'b001101000011: dataB <= 32'b00000100101101000010110010110000;
12'b001101000100: dataB <= 32'b00010001011010101110000111110111;
12'b001101000101: dataB <= 32'b00000101010010011111010110110110;
12'b001101000110: dataB <= 32'b01110010110110011001100010100100;
12'b001101000111: dataB <= 32'b00001110010010001010110111011010;
12'b001101001000: dataB <= 32'b10111011000111000010001110001011;
12'b001101001001: dataB <= 32'b00001101100101111100110110110011;
12'b001101001010: dataB <= 32'b11011001001111110011000001001000;
12'b001101001011: dataB <= 32'b00001111001011111010111010001100;
12'b001101001100: dataB <= 32'b10011100110001101101010101011110;
12'b001101001101: dataB <= 32'b00000010010110101101110011000011;
12'b001101001110: dataB <= 32'b01010100011111010001110110100100;
12'b001101001111: dataB <= 32'b00000100110100001001001111110011;
12'b001101010000: dataB <= 32'b10011110101101010101100111111000;
12'b001101010001: dataB <= 32'b00000011001001101010111101000000;
12'b001101010010: dataB <= 32'b00110110111101001100010111110010;
12'b001101010011: dataB <= 32'b00000111101101101000111100011010;
12'b001101010100: dataB <= 32'b01100001000011101010101000101010;
12'b001101010101: dataB <= 32'b00000111111001010011101101100011;
12'b001101010110: dataB <= 32'b01101011001011001011110100101100;
12'b001101010111: dataB <= 32'b00001010100110011010010110000100;
12'b001101011000: dataB <= 32'b00011001110001100010101011001110;
12'b001101011001: dataB <= 32'b00000101100001010010100001000110;
12'b001101011010: dataB <= 32'b11110010100110000000010111101000;
12'b001101011011: dataB <= 32'b00001011000010100100100110100001;
12'b001101011100: dataB <= 32'b00100000101101111001011011001010;
12'b001101011101: dataB <= 32'b00000101010110000101010111110100;
12'b001101011110: dataB <= 32'b01101001111010010100111011110110;
12'b001101011111: dataB <= 32'b00001000011110011001110010001111;
12'b001101100000: dataB <= 32'b10100101010110001000010110100110;
12'b001101100001: dataB <= 32'b00000101111110010001101001110100;
12'b001101100010: dataB <= 32'b11111100110010101101111100011011;
12'b001101100011: dataB <= 32'b00001000101011010110100111100001;
12'b001101100100: dataB <= 32'b10000011001111000101010010101100;
12'b001101100101: dataB <= 32'b00001000010101010101010000011100;
12'b001101100110: dataB <= 32'b10100000111110100010101011101110;
12'b001101100111: dataB <= 32'b00001111001100010100001010110011;
12'b001101101000: dataB <= 32'b11010000011110101110101000011001;
12'b001101101001: dataB <= 32'b00001101110101101111001101000000;
12'b001101101010: dataB <= 32'b01010000101101110000110011100011;
12'b001101101011: dataB <= 32'b00001111001011101110110001101011;
12'b001101101100: dataB <= 32'b00000111011111010001011110001011;
12'b001101101101: dataB <= 32'b00000111111000010011101111000111;
12'b001101101110: dataB <= 32'b10101001000001101010001101010010;
12'b001101101111: dataB <= 32'b00000010111001010011101111010100;
12'b001101110000: dataB <= 32'b01011001100010000000011101101111;
12'b001101110001: dataB <= 32'b00000001001000100111010010001110;
12'b001101110010: dataB <= 32'b00010010100110101101001000010011;
12'b001101110011: dataB <= 32'b00001100111010101011110111100100;
12'b001101110100: dataB <= 32'b00100011111000110101011000111010;
12'b001101110101: dataB <= 32'b00001100100100100100011001111110;
12'b001101110110: dataB <= 32'b11001111001110101000011010001010;
12'b001101110111: dataB <= 32'b00000010111010000101010101100100;
12'b001101111000: dataB <= 32'b01101101000101011000011001110000;
12'b001101111001: dataB <= 32'b00001101010111010111001010001011;
12'b001101111010: dataB <= 32'b11101111010110001000011001100111;
12'b001101111011: dataB <= 32'b00000011010110101001111001100011;
12'b001101111100: dataB <= 32'b00111101010101010001011110110001;
12'b001101111101: dataB <= 32'b00001011101111010100100101110011;
12'b001101111110: dataB <= 32'b10000110100010011101100000110010;
12'b001101111111: dataB <= 32'b00001011001011110100111010111100;
12'b001110000000: dataB <= 32'b11011111110010001001100110000110;
12'b001110000001: dataB <= 32'b00000010001111000011001110000101;
12'b001110000010: dataB <= 32'b11000011000111100011111011101111;
12'b001110000011: dataB <= 32'b00000110000111100110110100110100;
12'b001110000100: dataB <= 32'b01110011101010011110101011011101;
12'b001110000101: dataB <= 32'b00001111001110110100110001111101;
12'b001110000110: dataB <= 32'b01110100100110011100100111010001;
12'b001110000111: dataB <= 32'b00000100110011100001111011101010;
12'b001110001000: dataB <= 32'b11010010110011001110100000110000;
12'b001110001001: dataB <= 32'b00000101001011011010111100011001;
12'b001110001010: dataB <= 32'b01101001011010001101000010110000;
12'b001110001011: dataB <= 32'b00001001101000011100100011011110;
12'b001110001100: dataB <= 32'b00100001001010111010101000101100;
12'b001110001101: dataB <= 32'b00000101100001111101010111100101;
12'b001110001110: dataB <= 32'b01011100011101110100001101011000;
12'b001110001111: dataB <= 32'b00001100001110100110110111101010;
12'b001110010000: dataB <= 32'b01000101000101011101011000011000;
12'b001110010001: dataB <= 32'b00000111111110001001100010011110;
12'b001110010010: dataB <= 32'b10111101010111011010111011001010;
12'b001110010011: dataB <= 32'b00000100010111011001101001001010;
12'b001110010100: dataB <= 32'b11101101010000010010011101010111;
12'b001110010101: dataB <= 32'b00000110111110100111111001000010;
12'b001110010110: dataB <= 32'b11010001000001110100111011011101;
12'b001110010111: dataB <= 32'b00001010110101000010110010111101;
12'b001110011000: dataB <= 32'b11101110110010001000010101100001;
12'b001110011001: dataB <= 32'b00000100101100000100100111000000;
12'b001110011010: dataB <= 32'b01001111010010100110010111010111;
12'b001110011011: dataB <= 32'b00000100110001011101010010101110;
12'b001110011100: dataB <= 32'b11110010111110101001110100000011;
12'b001110011101: dataB <= 32'b00001101110101001010101111100010;
12'b001110011110: dataB <= 32'b00111001010011010010101110101110;
12'b001110011111: dataB <= 32'b00001110001000111100111110110100;
12'b001110100000: dataB <= 32'b00011001001011110011110010000110;
12'b001110100001: dataB <= 32'b00001111001110111011000110001101;
12'b001110100010: dataB <= 32'b00011110110001100101000100011100;
12'b001110100011: dataB <= 32'b00000001110100101001110111000100;
12'b001110100100: dataB <= 32'b00010110011011100010100111100100;
12'b001110100101: dataB <= 32'b00000100010010000111000111110100;
12'b001110100110: dataB <= 32'b01100000101101001101010110110111;
12'b001110100111: dataB <= 32'b00000011101000101011000001011000;
12'b001110101000: dataB <= 32'b01110111000101001011110111010010;
12'b001110101001: dataB <= 32'b00001000001101101001000000101001;
12'b001110101010: dataB <= 32'b01100001000011110011001001001010;
12'b001110101011: dataB <= 32'b00000110111000001111101001100011;
12'b001110101100: dataB <= 32'b01101001001111001100010101001010;
12'b001110101101: dataB <= 32'b00001011000111011110010110000100;
12'b001110101110: dataB <= 32'b10010011101101101010101011010000;
12'b001110101111: dataB <= 32'b00000110100001010110011100110101;
12'b001110110000: dataB <= 32'b00110100101110011000011000001000;
12'b001110110001: dataB <= 32'b00001100000011100110100110110010;
12'b001110110010: dataB <= 32'b11100000101110001001011011101011;
12'b001110110011: dataB <= 32'b00000100110100000101001011110100;
12'b001110110100: dataB <= 32'b01100011111010001101001011010111;
12'b001110110101: dataB <= 32'b00000110111110010101101101111111;
12'b001110110110: dataB <= 32'b10100011011010100000010111100110;
12'b001110110111: dataB <= 32'b00000100011101001101100001110100;
12'b001110111000: dataB <= 32'b10111100111110011110001011011100;
12'b001110111001: dataB <= 32'b00001001001011011010100011101010;
12'b001110111010: dataB <= 32'b11000011000010111101110011001010;
12'b001110111011: dataB <= 32'b00000111110101010011001100011011;
12'b001110111100: dataB <= 32'b00100000111110101010111011101111;
12'b001110111101: dataB <= 32'b00001111001111011010001010110100;
12'b001110111110: dataB <= 32'b01010100010110011110110111011001;
12'b001110111111: dataB <= 32'b00001101010111101101010101010000;
12'b001111000000: dataB <= 32'b01010010101010000000110101000010;
12'b001111000001: dataB <= 32'b00001111001101110000110101110011;
12'b001111000010: dataB <= 32'b01000011010011100001111110101101;
12'b001111000011: dataB <= 32'b00000111011000001111101010101111;
12'b001111000100: dataB <= 32'b00101001000001110010001100110100;
12'b001111000101: dataB <= 32'b00000001110110001111101011001101;
12'b001111000110: dataB <= 32'b01010111011110010000011101110001;
12'b001111000111: dataB <= 32'b00000010000110100101010010000110;
12'b001111001000: dataB <= 32'b11010100100010100101010111110011;
12'b001111001001: dataB <= 32'b00001011011100100101111011011100;
12'b001111001010: dataB <= 32'b00011101111000101100110111011010;
12'b001111001011: dataB <= 32'b00001101100110101000011101110110;
12'b001111001100: dataB <= 32'b11001101000110111000111010101011;
12'b001111001101: dataB <= 32'b00000001110111000011001001100100;
12'b001111001110: dataB <= 32'b01101011001001110000011001010001;
12'b001111001111: dataB <= 32'b00001100011001010111000110001011;
12'b001111010000: dataB <= 32'b10101101011010100000011010001000;
12'b001111010001: dataB <= 32'b00000010110100100011111001101011;
12'b001111010010: dataB <= 32'b00111001011101100001011110110100;
12'b001111010011: dataB <= 32'b00001011110000010110100001110011;
12'b001111010100: dataB <= 32'b11001010010110010101100000101111;
12'b001111010101: dataB <= 32'b00001011101101110101000110111100;
12'b001111010110: dataB <= 32'b11011001101110011001110111000101;
12'b001111010111: dataB <= 32'b00000010101101000011000001111101;
12'b001111011000: dataB <= 32'b01000010111011100100101011110000;
12'b001111011001: dataB <= 32'b00000111000110101000111000101100;
12'b001111011010: dataB <= 32'b01101101110010001110111010011110;
12'b001111011011: dataB <= 32'b00001111010001110110111001110101;
12'b001111011100: dataB <= 32'b00110110101110010100110110110000;
12'b001111011101: dataB <= 32'b00000100110010011011111011110011;
12'b001111011110: dataB <= 32'b01010100101110110111000000101101;
12'b001111011111: dataB <= 32'b00000101101010011010111100101001;
12'b001111100000: dataB <= 32'b11100101011110000101000010101110;
12'b001111100001: dataB <= 32'b00001010101001011110100011001110;
12'b001111100010: dataB <= 32'b10100001001011000011001000101100;
12'b001111100011: dataB <= 32'b00000111000001111001011111011101;
12'b001111100100: dataB <= 32'b00100000011101110100001100011010;
12'b001111100101: dataB <= 32'b00001100010000101000111011110011;
12'b001111100110: dataB <= 32'b10000100111101010101000111010111;
12'b001111100111: dataB <= 32'b00000110111110000111011010001110;
12'b001111101000: dataB <= 32'b01111001011111011011101011101011;
12'b001111101001: dataB <= 32'b00000011110101010101100101011010;
12'b001111101010: dataB <= 32'b10101011010100011001111100011001;
12'b001111101011: dataB <= 32'b00000101011110100001111001001010;
12'b001111101100: dataB <= 32'b00010000111101101100111010011110;
12'b001111101101: dataB <= 32'b00001010010101000100100110101110;
12'b001111101110: dataB <= 32'b01110000110110100000010111000001;
12'b001111101111: dataB <= 32'b00000101001011000110011111010001;
12'b001111110000: dataB <= 32'b10001111001110010110010110110110;
12'b001111110001: dataB <= 32'b00000100101111011011010010011110;
12'b001111110010: dataB <= 32'b01110011000110111010000101000001;
12'b001111110011: dataB <= 32'b00001101010111001100100111101011;
12'b001111110100: dataB <= 32'b01110111011011010011001110110000;
12'b001111110101: dataB <= 32'b00001111001010111101001010110100;
12'b001111110110: dataB <= 32'b00010111000111110100100011000100;
12'b001111110111: dataB <= 32'b00001111010001111011010010000101;
12'b001111111000: dataB <= 32'b01100000110001011101000010111010;
12'b001111111001: dataB <= 32'b00000001010010100011111011000100;
12'b001111111010: dataB <= 32'b10011010011011101011001000100100;
12'b001111111011: dataB <= 32'b00000100010001000110111111110100;
12'b001111111100: dataB <= 32'b01100000101101000101000110010111;
12'b001111111101: dataB <= 32'b00000100100110101011000101110000;
12'b001111111110: dataB <= 32'b11110111001101001011100111010010;
12'b001111111111: dataB <= 32'b00001000001101101001000000111000;
12'b010000000000: dataB <= 32'b00100001000011110011111001101011;
12'b010000000001: dataB <= 32'b00000101111000001011100001101011;
12'b010000000010: dataB <= 32'b01101001010011000100110101101010;
12'b010000000011: dataB <= 32'b00001100001000100010010110000100;
12'b010000000100: dataB <= 32'b00001111101001110010011011010001;
12'b010000000101: dataB <= 32'b00001000000001011000011100101101;
12'b010000000110: dataB <= 32'b01110110110110110000101001001000;
12'b010000000111: dataB <= 32'b00001101000101101000101010111010;
12'b010000001000: dataB <= 32'b10100010101110011001101100001101;
12'b010000001001: dataB <= 32'b00000100010011000011000011101101;
12'b010000001010: dataB <= 32'b01011101111010000101001010011000;
12'b010000001011: dataB <= 32'b00000101011110001111101001100111;
12'b010000001100: dataB <= 32'b01100001011010111000101000000110;
12'b010000001101: dataB <= 32'b00000011011011001001011001101100;
12'b010000001110: dataB <= 32'b01111101001010001110001001111101;
12'b010000001111: dataB <= 32'b00001001101100011100100011110011;
12'b010000010000: dataB <= 32'b01000010110110101110000011101000;
12'b010000010001: dataB <= 32'b00000111010101010001001000011011;
12'b010000010010: dataB <= 32'b01100000111110110011001011110001;
12'b010000010011: dataB <= 32'b00001111010010011110000110110100;
12'b010000010100: dataB <= 32'b01011000010010000111000110011000;
12'b010000010101: dataB <= 32'b00001100111001101011011001101000;
12'b010000010110: dataB <= 32'b01010100100110011001000110100001;
12'b010000010111: dataB <= 32'b00001111010000110000111101110011;
12'b010000011000: dataB <= 32'b10000011001011101010011110110000;
12'b010000011001: dataB <= 32'b00000110011000001011100010010111;
12'b010000011010: dataB <= 32'b01101001000110000010001100010101;
12'b010000011011: dataB <= 32'b00000001010100001011100011000101;
12'b010000011100: dataB <= 32'b01010011011010101000101101010011;
12'b010000011101: dataB <= 32'b00000011000100100011010101110110;
12'b010000011110: dataB <= 32'b01010110011110011101100111010011;
12'b010000011111: dataB <= 32'b00001010011101011111111011010101;
12'b010000100000: dataB <= 32'b00010111111000101100010110011010;
12'b010000100001: dataB <= 32'b00001110101000101100100001100110;
12'b010000100010: dataB <= 32'b10001100111111010001011011001100;
12'b010000100011: dataB <= 32'b00000000110101000010111101011100;
12'b010000100100: dataB <= 32'b10101011001110001000011001010001;
12'b010000100101: dataB <= 32'b00001011011011010111000010010011;
12'b010000100110: dataB <= 32'b10101001011110111000101011001001;
12'b010000100111: dataB <= 32'b00000010110010011101111001101011;
12'b010000101000: dataB <= 32'b00110101101001110001001110010110;
12'b010000101001: dataB <= 32'b00001011010010011010011101111011;
12'b010000101010: dataB <= 32'b00001110001110000101110000101100;
12'b010000101011: dataB <= 32'b00001011101110110101001110110101;
12'b010000101100: dataB <= 32'b10010101101010101001111000000101;
12'b010000101101: dataB <= 32'b00000010101011000010110101101101;
12'b010000101110: dataB <= 32'b11000010101111011101001011010010;
12'b010000101111: dataB <= 32'b00001000000110101000111100101011;
12'b010000110000: dataB <= 32'b00101001110101110110111000111110;
12'b010000110001: dataB <= 32'b00001111010100110111000101101101;
12'b010000110010: dataB <= 32'b11111000110110001100110110110000;
12'b010000110011: dataB <= 32'b00000100010000010101111011110011;
12'b010000110100: dataB <= 32'b11010110101010100111010000101010;
12'b010000110101: dataB <= 32'b00000110001001011010111101000000;
12'b010000110110: dataB <= 32'b01100011011101111101000011001100;
12'b010000110111: dataB <= 32'b00001011001010100010100010111111;
12'b010000111000: dataB <= 32'b00011111001011000011101001001100;
12'b010000111001: dataB <= 32'b00001000100001110101101011001110;
12'b010000111010: dataB <= 32'b11100100011101110011111010111011;
12'b010000111011: dataB <= 32'b00001100010010101000111111110011;
12'b010000111100: dataB <= 32'b10000100110001001100110110110111;
12'b010000111101: dataB <= 32'b00000101011101000101001101111110;
12'b010000111110: dataB <= 32'b00110101101011100100001100001101;
12'b010000111111: dataB <= 32'b00000011010100010001100001100010;
12'b010001000000: dataB <= 32'b01101001011000101001011011011011;
12'b010001000001: dataB <= 32'b00000100011100011011111001010010;
12'b010001000010: dataB <= 32'b01010010110101100100101000111110;
12'b010001000011: dataB <= 32'b00001001010110000110011110100110;
12'b010001000100: dataB <= 32'b00110000111110111000101000100001;
12'b010001000101: dataB <= 32'b00000101101010001010010111100010;
12'b010001000110: dataB <= 32'b10001101000110000110010101110101;
12'b010001000111: dataB <= 32'b00000100101110011001001110001110;
12'b010001001000: dataB <= 32'b00110001001111000010100110100001;
12'b010001001001: dataB <= 32'b00001100111001010000100011101100;
12'b010001001010: dataB <= 32'b10110011100011011011101110110011;
12'b010001001011: dataB <= 32'b00001111001101111011010110110100;
12'b010001001100: dataB <= 32'b00010111000011110101000100000010;
12'b010001001101: dataB <= 32'b00001111010100111001011001111101;
12'b010001001110: dataB <= 32'b11100010110001010100110001111000;
12'b010001001111: dataB <= 32'b00000001001111011101111011000100;
12'b010001010000: dataB <= 32'b01011110011011101011111001100101;
12'b010001010001: dataB <= 32'b00000100001111001000110011101101;
12'b010001010010: dataB <= 32'b01100010101100111100100101110110;
12'b010001010011: dataB <= 32'b00000101100101101001001010001000;
12'b010001010100: dataB <= 32'b10110101010101001011010110110001;
12'b010001010101: dataB <= 32'b00001000001101101001000101001000;
12'b010001010110: dataB <= 32'b00100001000011110100101010001100;
12'b010001010111: dataB <= 32'b00000101010111001001010101110011;
12'b010001011000: dataB <= 32'b01100111010111000101010110101001;
12'b010001011001: dataB <= 32'b00001100101010100110011001111100;
12'b010001011010: dataB <= 32'b10001011100001111010011011010010;
12'b010001011011: dataB <= 32'b00001001100001011100011000101100;
12'b010001011100: dataB <= 32'b11110110111111000000111001101001;
12'b010001011101: dataB <= 32'b00001110001000101010101111000010;
12'b010001011110: dataB <= 32'b00100100110010101001111100001110;
12'b010001011111: dataB <= 32'b00000100010010000100110111100110;
12'b010001100000: dataB <= 32'b00010111111010000101001001011001;
12'b010001100001: dataB <= 32'b00000100011100001011100001010111;
12'b010001100010: dataB <= 32'b01011101011011001001001001000110;
12'b010001100011: dataB <= 32'b00000010011001000111010001101100;
12'b010001100100: dataB <= 32'b11111011010110000110001000011110;
12'b010001100101: dataB <= 32'b00001001101100100000011111110011;
12'b010001100110: dataB <= 32'b10000010101010011110010100100111;
12'b010001100111: dataB <= 32'b00000110110101010001000000100010;
12'b010001101000: dataB <= 32'b10100000111110110011011011110010;
12'b010001101001: dataB <= 32'b00001110110101100100001010101100;
12'b010001101010: dataB <= 32'b01011100010001110111000101111000;
12'b010001101011: dataB <= 32'b00001011111010100111011110000000;
12'b010001101100: dataB <= 32'b00010110100010101001010111100001;
12'b010001101101: dataB <= 32'b00001111010011110001000101111011;
12'b010001101110: dataB <= 32'b10000010111111110011001110110011;
12'b010001101111: dataB <= 32'b00000101010111001001011010000111;
12'b010001110000: dataB <= 32'b11100111001010001010001011110111;
12'b010001110001: dataB <= 32'b00000001010001001001011010111101;
12'b010001110010: dataB <= 32'b00010001010111000000111101010101;
12'b010001110011: dataB <= 32'b00000100000010100001010101100110;
12'b010001110100: dataB <= 32'b11011010011110010101100111010011;
12'b010001110101: dataB <= 32'b00001000111101011001111011001101;
12'b010001110110: dataB <= 32'b11010001110100101011100101011001;
12'b010001110111: dataB <= 32'b00001111001011101110100101010101;
12'b010001111000: dataB <= 32'b01001100111011100001111011001101;
12'b010001111001: dataB <= 32'b00000000110010000010110001011100;
12'b010001111010: dataB <= 32'b10101001010010100000011001010010;
12'b010001111011: dataB <= 32'b00001010011100010110111110010011;
12'b010001111100: dataB <= 32'b01100111100011001001001011101010;
12'b010001111101: dataB <= 32'b00000010010000010111111001101011;
12'b010001111110: dataB <= 32'b00110001110010000001001101011001;
12'b010001111111: dataB <= 32'b00001011010011011100011110000011;
12'b010010000000: dataB <= 32'b10010010001001111101110001001001;
12'b010010000001: dataB <= 32'b00001100010000110011010110101101;
12'b010010000010: dataB <= 32'b10010001100110110010011001000101;
12'b010010000011: dataB <= 32'b00000011001001000010101101100101;
12'b010010000100: dataB <= 32'b01000100100011010101101011010011;
12'b010010000101: dataB <= 32'b00001000100110101000111100101011;
12'b010010000110: dataB <= 32'b00100011110101100110100111011110;
12'b010010000111: dataB <= 32'b00001110110110110101001101100101;
12'b010010001000: dataB <= 32'b10111001000010001100110110110000;
12'b010010001001: dataB <= 32'b00000100001111010001110011110100;
12'b010010001010: dataB <= 32'b01011000100110001111010001101000;
12'b010010001011: dataB <= 32'b00000110101001011100111001010000;
12'b010010001100: dataB <= 32'b10011111100001110101000011101010;
12'b010010001101: dataB <= 32'b00001011101100100100100010100111;
12'b010010001110: dataB <= 32'b10011111001011000011111001101101;
12'b010010001111: dataB <= 32'b00001010000001110001110010111110;
12'b010010010000: dataB <= 32'b10100110100001110011111001111100;
12'b010010010001: dataB <= 32'b00001011110011101000111111110100;
12'b010010010010: dataB <= 32'b10000110101001001100100101110110;
12'b010010010011: dataB <= 32'b00000011111100000011000001101110;
12'b010010010100: dataB <= 32'b00110001110011011100101100001110;
12'b010010010101: dataB <= 32'b00000010110010001111011001101010;
12'b010010010110: dataB <= 32'b00100101011101000000111010011100;
12'b010010010111: dataB <= 32'b00000010111010010101110101011010;
12'b010010011000: dataB <= 32'b10010010110001100100010111011110;
12'b010010011001: dataB <= 32'b00001000110111001010010110010110;
12'b010010011010: dataB <= 32'b10110001000111001001001010000001;
12'b010010011011: dataB <= 32'b00000110001001010000001111110010;
12'b010010011100: dataB <= 32'b10001100111101110110010101010101;
12'b010010011101: dataB <= 32'b00000101001101011001001101110110;
12'b010010011110: dataB <= 32'b11110001010011001011001000000001;
12'b010010011111: dataB <= 32'b00001011111010010010011011101100;
12'b010010100000: dataB <= 32'b11101111101011011100001110010101;
12'b010010100001: dataB <= 32'b00001111010000111001100010101100;
12'b010010100010: dataB <= 32'b00010111000011100101110101100001;
12'b010010100011: dataB <= 32'b00001110110111110101100101110101;
12'b010010100100: dataB <= 32'b01100010110001010100010001010110;
12'b010010100101: dataB <= 32'b00000001001100010111110110111101;
12'b010010100110: dataB <= 32'b00100010011011101100011010100101;
12'b010010100111: dataB <= 32'b00000100001110001010101011100110;
12'b010010101000: dataB <= 32'b01100100110000111100010100110101;
12'b010010101001: dataB <= 32'b00000110100100101001001110100000;
12'b010010101010: dataB <= 32'b01110001011101010011000110110001;
12'b010010101011: dataB <= 32'b00001000101110100111001001100000;
12'b010010101100: dataB <= 32'b00100001000011101101011010101101;
12'b010010101101: dataB <= 32'b00000100110110000111001101110011;
12'b010010101110: dataB <= 32'b01100011010110110101100111001000;
12'b010010101111: dataB <= 32'b00001101001100101010011101111100;
12'b010010110000: dataB <= 32'b00001001011010001010011010110011;
12'b010010110001: dataB <= 32'b00001011000010100000011000100100;
12'b010010110010: dataB <= 32'b01110111000111010001011010001010;
12'b010010110011: dataB <= 32'b00001111001010101100110011001011;
12'b010010110100: dataB <= 32'b11100110110010111010001100010000;
12'b010010110101: dataB <= 32'b00000011110000000100101011010110;
12'b010010110110: dataB <= 32'b10010001110101111101001000011010;
12'b010010110111: dataB <= 32'b00000010111011001001011000111110;
12'b010010111000: dataB <= 32'b00011011010111011001101010000111;
12'b010010111001: dataB <= 32'b00000001010111000101000101101100;
12'b010010111010: dataB <= 32'b10111001100001110110000111011110;
12'b010010111011: dataB <= 32'b00001010001101100010100011110100;
12'b010010111100: dataB <= 32'b00000110100010001110010101000110;
12'b010010111101: dataB <= 32'b00000110010100010000111100101010;
12'b010010111110: dataB <= 32'b11100000111110110011101011010100;
12'b010010111111: dataB <= 32'b00001110011000101010001010101100;
12'b010011000000: dataB <= 32'b01100000010001100110110100110111;
12'b010011000001: dataB <= 32'b00001010011100100101011110011000;
12'b010011000010: dataB <= 32'b00011010011110111001101001000001;
12'b010011000011: dataB <= 32'b00001110110110110001001010000011;
12'b010011000100: dataB <= 32'b10000010110011110011111110010101;
12'b010011000101: dataB <= 32'b00000100110110000111001101101111;
12'b010011000110: dataB <= 32'b00100111001110011010001010111000;
12'b010011000111: dataB <= 32'b00000001001110000111001110101110;
12'b010011001000: dataB <= 32'b11001111001111010001011100010111;
12'b010011001001: dataB <= 32'b00000101100001011111010101011101;
12'b010011001010: dataB <= 32'b01011110011010001101100110110010;
12'b010011001011: dataB <= 32'b00000111011101010101110110111110;
12'b010011001100: dataB <= 32'b10001101101100101011000100111000;
12'b010011001101: dataB <= 32'b00001111001110110000101101001101;
12'b010011001110: dataB <= 32'b00001110110011101010011011001110;
12'b010011001111: dataB <= 32'b00000000101111000100101001010100;
12'b010011010000: dataB <= 32'b11100111010110111000101000110010;
12'b010011010001: dataB <= 32'b00001000111101010110111010010011;
12'b010011010010: dataB <= 32'b01100011100011011001101100001100;
12'b010011010011: dataB <= 32'b00000010001110010001110101110011;
12'b010011010100: dataB <= 32'b00101101110110010001001100011010;
12'b010011010101: dataB <= 32'b00001010110100100000011110001011;
12'b010011010110: dataB <= 32'b11011000000101101101100010000110;
12'b010011010111: dataB <= 32'b00001011110001110001011010100101;
12'b010011011000: dataB <= 32'b01001101011110111010101010000110;
12'b010011011001: dataB <= 32'b00000100000111000110100001011101;
12'b010011011010: dataB <= 32'b11001000011011000110001010110100;
12'b010011011011: dataB <= 32'b00001001100111101001000000110010;
12'b010011011100: dataB <= 32'b11011101110101010110010101111110;
12'b010011011101: dataB <= 32'b00001101111001110011010101011100;
12'b010011011110: dataB <= 32'b00111001001010000101000110101111;
12'b010011011111: dataB <= 32'b00000100101101001011101111110101;
12'b010011100000: dataB <= 32'b01011010100101110111010010000101;
12'b010011100001: dataB <= 32'b00000111001001011100111001101000;
12'b010011100010: dataB <= 32'b10011101011101110100110100001000;
12'b010011100011: dataB <= 32'b00001011101101101000100110001111;
12'b010011100100: dataB <= 32'b11011101001011000100011001101101;
12'b010011100101: dataB <= 32'b00001011100010101101110110101110;
12'b010011100110: dataB <= 32'b00101010100101110011111000011101;
12'b010011100111: dataB <= 32'b00001011010101101001000011110101;
12'b010011101000: dataB <= 32'b01001010011101001100010101010101;
12'b010011101001: dataB <= 32'b00000010111010000010111001011110;
12'b010011101010: dataB <= 32'b11101101110111010101011100010000;
12'b010011101011: dataB <= 32'b00000010110000001101010101111001;
12'b010011101100: dataB <= 32'b11100011011101010000011000111101;
12'b010011101101: dataB <= 32'b00000001111000001111110001101001;
12'b010011101110: dataB <= 32'b10010100101101100100010101111110;
12'b010011101111: dataB <= 32'b00001000010111010000001110000110;
12'b010011110000: dataB <= 32'b01110001001011011001101011100010;
12'b010011110001: dataB <= 32'b00000110101001010100000111110011;
12'b010011110010: dataB <= 32'b10001100110101100110010100110011;
12'b010011110011: dataB <= 32'b00000101001100010111001001100110;
12'b010011110100: dataB <= 32'b01101111011011001011101001100001;
12'b010011110101: dataB <= 32'b00001010011100010110010111100101;
12'b010011110110: dataB <= 32'b00101011101111011100101101011000;
12'b010011110111: dataB <= 32'b00001111010011110101101010100101;
12'b010011111000: dataB <= 32'b11010110111111011110010111000001;
12'b010011111001: dataB <= 32'b00001101111001110001101001110100;
12'b010011111010: dataB <= 32'b10100100110101001100000000110011;
12'b010011111011: dataB <= 32'b00000001101010010011110010110101;
12'b010011111100: dataB <= 32'b10100110011011100101001011100111;
12'b010011111101: dataB <= 32'b00000100001100001100100011010110;
12'b010011111110: dataB <= 32'b10100110110000111011110100010100;
12'b010011111111: dataB <= 32'b00000111100100100111010010111000;
12'b010100000000: dataB <= 32'b01101111100101011010110110110000;
12'b010100000001: dataB <= 32'b00001000101110100111001101111000;
12'b010100000010: dataB <= 32'b11100001000011100110001010101110;
12'b010100000011: dataB <= 32'b00000011110100000101000001111010;
12'b010100000100: dataB <= 32'b01100001011010101101110111101000;
12'b010100000101: dataB <= 32'b00001101101110101110100001111100;
12'b010100000110: dataB <= 32'b10000111001110010010101010010100;
12'b010100000111: dataB <= 32'b00001100100100100100011000100011;
12'b010100001000: dataB <= 32'b11110101010011100010001010101011;
12'b010100001001: dataB <= 32'b00001111001101101100110111010011;
12'b010100001010: dataB <= 32'b00100110110111000010101100010010;
12'b010100001011: dataB <= 32'b00000011101110001000100010111111;
12'b010100001100: dataB <= 32'b01001101101101110101000111011010;
12'b010100001101: dataB <= 32'b00000001111000000111010000101110;
12'b010100001110: dataB <= 32'b00011001010111101010011011001000;
12'b010100001111: dataB <= 32'b00000000110100000100111101101100;
12'b010100010000: dataB <= 32'b01110101101001100110000101111101;
12'b010100010001: dataB <= 32'b00001010001110100110100011101101;
12'b010100010010: dataB <= 32'b10001010010101111110100110000101;
12'b010100010011: dataB <= 32'b00000101110011010000110100111001;
12'b010100010100: dataB <= 32'b00100000111110111100001010110101;
12'b010100010101: dataB <= 32'b00001101011010101110010010100101;
12'b010100010110: dataB <= 32'b10100100010001010110100100010101;
12'b010100010111: dataB <= 32'b00001001011100100001011110110000;
12'b010100011000: dataB <= 32'b00011110011111001010001010100010;
12'b010100011001: dataB <= 32'b00001101111000101111010010000011;
12'b010100011010: dataB <= 32'b01000100100111110100101101010111;
12'b010100011011: dataB <= 32'b00000100010100000111000101010111;
12'b010100011100: dataB <= 32'b01100101001110100010011001111001;
12'b010100011101: dataB <= 32'b00000001001100000111000110011110;
12'b010100011110: dataB <= 32'b10001111000111100001111011011001;
12'b010100011111: dataB <= 32'b00000111000001011101010101001101;
12'b010100100000: dataB <= 32'b10100010011001111101110110110010;
12'b010100100001: dataB <= 32'b00000110011101001111110010110110;
12'b010100100010: dataB <= 32'b00001001100100110010100011110110;
12'b010100100011: dataB <= 32'b00001111010001110010110101000101;
12'b010100100100: dataB <= 32'b11010000101011110011001011110000;
12'b010100100101: dataB <= 32'b00000000101100000110011101010011;
12'b010100100110: dataB <= 32'b11100101010111001001001000110010;
12'b010100100111: dataB <= 32'b00000111111101010110110110010011;
12'b010100101000: dataB <= 32'b01011111100111101010011100001110;
12'b010100101001: dataB <= 32'b00000010101100001101101101110011;
12'b010100101010: dataB <= 32'b00100111111010100001011011011100;
12'b010100101011: dataB <= 32'b00001010010101100100011110001011;
12'b010100101100: dataB <= 32'b11011110000101100101100010100100;
12'b010100101101: dataB <= 32'b00001011110011101101100010010101;
12'b010100101110: dataB <= 32'b00001011011011000011001011000111;
12'b010100101111: dataB <= 32'b00000101000110001000011001010101;
12'b010100110000: dataB <= 32'b01001100010010111110101010010101;
12'b010100110001: dataB <= 32'b00001010101000101001000100111010;
12'b010100110010: dataB <= 32'b10011001110101000110000100011101;
12'b010100110011: dataB <= 32'b00001100111011110001011101011100;
12'b010100110100: dataB <= 32'b11110111010001111101000110101111;
12'b010100110101: dataB <= 32'b00000100101100000111100011100101;
12'b010100110110: dataB <= 32'b01011110100101100111010011100011;
12'b010100110111: dataB <= 32'b00001000001000011100111010000000;
12'b010100111000: dataB <= 32'b10011001011101101100110101000111;
12'b010100111001: dataB <= 32'b00001011101111101010101001110111;
12'b010100111010: dataB <= 32'b00011101001011000100111001101110;
12'b010100111011: dataB <= 32'b00001100100100100111111010011111;
12'b010100111100: dataB <= 32'b11101100101001110011110111011101;
12'b010100111101: dataB <= 32'b00001010110110101001000111100101;
12'b010100111110: dataB <= 32'b00001100010101000011110100110100;
12'b010100111111: dataB <= 32'b00000001111000000100101101001110;
12'b010101000000: dataB <= 32'b11100111111011001101111100010010;
12'b010101000001: dataB <= 32'b00000010101101001011001110001001;
12'b010101000010: dataB <= 32'b11011111100001101000010111111101;
12'b010101000011: dataB <= 32'b00000001010110001011101001111001;
12'b010101000100: dataB <= 32'b10010110101001100100000100011101;
12'b010101000101: dataB <= 32'b00000111010111010100000101101110;
12'b010101000110: dataB <= 32'b00101111010011101010011100100100;
12'b010101000111: dataB <= 32'b00000111101001011010000111110100;
12'b010101001000: dataB <= 32'b01001110101101010110000100110010;
12'b010101001001: dataB <= 32'b00000101101011010111000101010110;
12'b010101001010: dataB <= 32'b11101011011111010100001011000010;
12'b010101001011: dataB <= 32'b00001001011100011010010111010101;
12'b010101001100: dataB <= 32'b01100111110011010101001100111010;
12'b010101001101: dataB <= 32'b00001110110110110001110010011101;
12'b010101001110: dataB <= 32'b11010110111011001110111000100001;
12'b010101001111: dataB <= 32'b00001100111011101101110001101100;
12'b010101010000: dataB <= 32'b11100100110101001011110000110000;
12'b010101010001: dataB <= 32'b00000010101000001111101010100101;
12'b010101010010: dataB <= 32'b00101010011111011101101100101001;
12'b010101010011: dataB <= 32'b00000100101011010000011011000111;
12'b010101010100: dataB <= 32'b00100110110100111011010100010010;
12'b010101010101: dataB <= 32'b00001000100100100101010011001001;
12'b010101010110: dataB <= 32'b01101011101001100010100110110000;
12'b010101010111: dataB <= 32'b00001000101110100101001110010000;
12'b010101011000: dataB <= 32'b11100001000011010110101010101111;
12'b010101011001: dataB <= 32'b00000011110010000100111010000010;
12'b010101011010: dataB <= 32'b01011111011010011110001000101000;
12'b010101011011: dataB <= 32'b00001101110000110000101001111100;
12'b010101011100: dataB <= 32'b00000111000110011010101001110101;
12'b010101011101: dataB <= 32'b00001101100101101000011100101011;
12'b010101011110: dataB <= 32'b01110011011011110010101011001100;
12'b010101011111: dataB <= 32'b00001111010000101100111111010100;
12'b010101100000: dataB <= 32'b00011010110001010001111001000111;
12'b010101100001: dataB <= 32'b00000111011000010001101111100010;
12'b010101100010: dataB <= 32'b10110111100110100100011101010001;
12'b010101100011: dataB <= 32'b00001100011100101001110011001110;
12'b010101100100: dataB <= 32'b10101011001101001000100100001001;
12'b010101100101: dataB <= 32'b00001010011110011111110110000100;
12'b010101100110: dataB <= 32'b10110100010111000100111110110100;
12'b010101100111: dataB <= 32'b00000111001011010000110010101000;
12'b010101101000: dataB <= 32'b00001011101011010100000010110011;
12'b010101101001: dataB <= 32'b00001001110100011011011100110110;
12'b010101101010: dataB <= 32'b11011110111110000010001010101010;
12'b010101101011: dataB <= 32'b00001101000101001000100010100010;
12'b010101101100: dataB <= 32'b01001000110111010101011010110111;
12'b010101101101: dataB <= 32'b00001110001101101110111100010010;
12'b010101101110: dataB <= 32'b11001111000001000001100001001010;
12'b010101101111: dataB <= 32'b00001100000100101000100001100011;
12'b010101110000: dataB <= 32'b01010011110110010000011011100101;
12'b010101110001: dataB <= 32'b00001010010111100011110011101101;
12'b010101110010: dataB <= 32'b00100110110101001010111100101100;
12'b010101110011: dataB <= 32'b00000110011101100011110011001011;
12'b010101110100: dataB <= 32'b10100011100000111000111100101001;
12'b010101110101: dataB <= 32'b00000000110001101011000110110101;
12'b010101110110: dataB <= 32'b01001100111010111100001001010010;
12'b010101110111: dataB <= 32'b00001110110011111001100011010010;
12'b010101111000: dataB <= 32'b11110011101101010110011011011000;
12'b010101111001: dataB <= 32'b00001000100001011010011010100101;
12'b010101111010: dataB <= 32'b01010101011101100000011000001000;
12'b010101111011: dataB <= 32'b00000110011110001111110001111101;
12'b010101111100: dataB <= 32'b01101010110100100001101001001110;
12'b010101111101: dataB <= 32'b00001110110000011011010001111011;
12'b010101111110: dataB <= 32'b01110011000001001000100111000111;
12'b010101111111: dataB <= 32'b00000110011010110111100101101100;
12'b010110000000: dataB <= 32'b10111100110000101010111110001001;
12'b010110000001: dataB <= 32'b00001010101011001110110101100011;
12'b010110000010: dataB <= 32'b01000011000010110100110010011010;
12'b010110000011: dataB <= 32'b00001001101000110000100110111011;
12'b010110000100: dataB <= 32'b01101101101001100001110011101001;
12'b010110000101: dataB <= 32'b00000011010101001101101110100101;
12'b010110000110: dataB <= 32'b00001001100111010010001010101011;
12'b010110000111: dataB <= 32'b00000100001010100010101101001110;
12'b010110001000: dataB <= 32'b00111011001111000101111110110111;
12'b010110001001: dataB <= 32'b00001101100110101110011110010101;
12'b010110001010: dataB <= 32'b11101000010010100100000111110010;
12'b010110001011: dataB <= 32'b00000110010110110001110010111000;
12'b010110001100: dataB <= 32'b11010011000011101100110001111000;
12'b010110001101: dataB <= 32'b00000100001111011101000100001011;
12'b010110001110: dataB <= 32'b01101111001110011100100011110101;
12'b010110001111: dataB <= 32'b00000111101000010100101011110100;
12'b010110010000: dataB <= 32'b00100101000110011001110111001100;
12'b010110010001: dataB <= 32'b00000010000110111100110011100011;
12'b010110010010: dataB <= 32'b11010100100101111100011110110001;
12'b010110010011: dataB <= 32'b00001011001010100010101110111000;
12'b010110010100: dataB <= 32'b10001011100101111101111010010110;
12'b010110010101: dataB <= 32'b00001100011100010111110111000101;
12'b010110010110: dataB <= 32'b10111100110010111001101001000111;
12'b010110010111: dataB <= 32'b00000110111010100111101000111011;
12'b010110011000: dataB <= 32'b00110001000000001100101110110000;
12'b010110011001: dataB <= 32'b00001011011101110101101000111100;
12'b010110011010: dataB <= 32'b10010101010010000100111110110111;
12'b010110011011: dataB <= 32'b00001011110001000011010111010100;
12'b010110011100: dataB <= 32'b01101000100001001000100010000110;
12'b010110011101: dataB <= 32'b00000100110000000011001010000000;
12'b010110011110: dataB <= 32'b01010111100011000101011001010110;
12'b010110011111: dataB <= 32'b00000101110100100011010011001101;
12'b010110100000: dataB <= 32'b01101110101010000001010001001001;
12'b010110100001: dataB <= 32'b00001110001101001011001010111001;
12'b010110100010: dataB <= 32'b00111000110010100001011101000110;
12'b010110100011: dataB <= 32'b00001011000010111000011110101011;
12'b010110100100: dataB <= 32'b10011101010011011001100000101110;
12'b010110100101: dataB <= 32'b00001101100110111000100110011100;
12'b010110100110: dataB <= 32'b11011010110101111101101000011110;
12'b010110100111: dataB <= 32'b00000100011010110101100010111010;
12'b010110101000: dataB <= 32'b11001110101010110001000100100110;
12'b010110101001: dataB <= 32'b00000101110110001101011111100001;
12'b010110101010: dataB <= 32'b10011010110001101110001001010111;
12'b010110101011: dataB <= 32'b00000010001110101000110100100001;
12'b010110101100: dataB <= 32'b01110100101001010100111000010010;
12'b010110101101: dataB <= 32'b00000111001110100110110100001011;
12'b010110101110: dataB <= 32'b11100000111111010001010111101010;
12'b010110101111: dataB <= 32'b00001001011000011101110101011011;
12'b010110110000: dataB <= 32'b00101101000011000011000100001110;
12'b010110110001: dataB <= 32'b00001000000100010100011110001100;
12'b010110110010: dataB <= 32'b10100011110001010011001010101100;
12'b010110110011: dataB <= 32'b00000010100100001110101101100110;
12'b010110110100: dataB <= 32'b01101100011001010000010110001001;
12'b010110110101: dataB <= 32'b00001000000001011110100110001001;
12'b010110110110: dataB <= 32'b01011000110001000010001000000111;
12'b010110110111: dataB <= 32'b00001000011000010101110111011001;
12'b010110111000: dataB <= 32'b00111011011110100100001101001111;
12'b010110111001: dataB <= 32'b00001101111010101101101111010110;
12'b010110111010: dataB <= 32'b10101011001000110001000011101011;
12'b010110111011: dataB <= 32'b00001011111101100011110110000100;
12'b010110111100: dataB <= 32'b01110000001111000100011111010001;
12'b010110111101: dataB <= 32'b00000110101011010000111010010000;
12'b010110111110: dataB <= 32'b10010001110011001011100011010101;
12'b010110111111: dataB <= 32'b00001010010011011111011101000110;
12'b010111000000: dataB <= 32'b10011110111101110010011010001001;
12'b010111000001: dataB <= 32'b00001100000011000100101010011010;
12'b010111000010: dataB <= 32'b00001000111111011100111011110110;
12'b010111000011: dataB <= 32'b00001110001011101110110100001011;
12'b010111000100: dataB <= 32'b11001111001000110010000000101101;
12'b010111000101: dataB <= 32'b00001011000010100100011101100011;
12'b010111000110: dataB <= 32'b10011001111001111000011010100011;
12'b010111000111: dataB <= 32'b00001011010110100111110011110100;
12'b010111001000: dataB <= 32'b10100110110001000011001100001010;
12'b010111001001: dataB <= 32'b00000111011101100111110011000010;
12'b010111001010: dataB <= 32'b00100111100000101001011011100111;
12'b010111001011: dataB <= 32'b00000000110100101011000010111101;
12'b010111001100: dataB <= 32'b00001101000010110011101001010010;
12'b010111001101: dataB <= 32'b00001110110001111011010111001010;
12'b010111001110: dataB <= 32'b10110111100101100110101100010110;
12'b010111001111: dataB <= 32'b00000111000001010110011110110101;
12'b010111010000: dataB <= 32'b01011001100001001000100111001001;
12'b010111010001: dataB <= 32'b00000111111110010101110110000101;
12'b010111010010: dataB <= 32'b01101010110000010010001001001110;
12'b010111010011: dataB <= 32'b00001110101110011101010001111011;
12'b010111010100: dataB <= 32'b01110000111000110001000110000111;
12'b010111010101: dataB <= 32'b00000111011011111011011101101100;
12'b010111010110: dataB <= 32'b10111010100100100011011101000111;
12'b010111010111: dataB <= 32'b00001010001010001110111101100011;
12'b010111011000: dataB <= 32'b11000011001110110100100011011011;
12'b010111011001: dataB <= 32'b00001000101000101100011110111010;
12'b010111011010: dataB <= 32'b00101111100101010010000011001011;
12'b010111011011: dataB <= 32'b00000011110111010001110010101101;
12'b010111011100: dataB <= 32'b01001101101111000001111010001010;
12'b010111011101: dataB <= 32'b00000011101100100000101101011110;
12'b010111011110: dataB <= 32'b00111011000111001101011111010100;
12'b010111011111: dataB <= 32'b00001100100100101010011010011101;
12'b010111100000: dataB <= 32'b01100100001110100011110111110010;
12'b010111100001: dataB <= 32'b00000110110110110111101010100000;
12'b010111100010: dataB <= 32'b10010011001011101100010010111011;
12'b010111100011: dataB <= 32'b00000100110001011101000100001100;
12'b010111100100: dataB <= 32'b10101111000110011100010100010111;
12'b010111100101: dataB <= 32'b00000110101000010010101111110011;
12'b010111100110: dataB <= 32'b10100101000110001001110110101100;
12'b010111100111: dataB <= 32'b00000001001000111010100111011010;
12'b010111101000: dataB <= 32'b01010010101001111100011110101111;
12'b010111101001: dataB <= 32'b00001010101001100000101110100000;
12'b010111101010: dataB <= 32'b00001111101010001101101010110101;
12'b010111101011: dataB <= 32'b00001101011010011101111011001101;
12'b010111101100: dataB <= 32'b00111010100110101001011000000111;
12'b010111101101: dataB <= 32'b00001000011010101011100100111100;
12'b010111101110: dataB <= 32'b10101110111000001101011110101110;
12'b010111101111: dataB <= 32'b00001100011100111001100000111100;
12'b010111110000: dataB <= 32'b11010111010110001100111111010100;
12'b010111110001: dataB <= 32'b00001011101111000111011111010011;
12'b010111110010: dataB <= 32'b01100100011100110001000001001000;
12'b010111110011: dataB <= 32'b00000100110010000011010101101000;
12'b010111110100: dataB <= 32'b11011011100111001100111001110110;
12'b010111110101: dataB <= 32'b00000110010101100101010011010100;
12'b010111110110: dataB <= 32'b11101100100001110001100000101100;
12'b010111110111: dataB <= 32'b00001110001011001011010010101000;
12'b010111111000: dataB <= 32'b11110110101010010001001100000101;
12'b010111111001: dataB <= 32'b00001001100001110100010110100010;
12'b010111111010: dataB <= 32'b01011111010011001001000000110001;
12'b010111111011: dataB <= 32'b00001100100100110100011110011100;
12'b010111111100: dataB <= 32'b01011010110110000101101001111110;
12'b010111111101: dataB <= 32'b00000101011100111001011010110010;
12'b010111111110: dataB <= 32'b01001100110010100000110011101000;
12'b010111111111: dataB <= 32'b00000110010111010001100111010001;
12'b011000000000: dataB <= 32'b00011000110001111110001010010111;
12'b011000000001: dataB <= 32'b00000010010000101000110000010010;
12'b011000000010: dataB <= 32'b00110010100001011101001000010010;
12'b011000000011: dataB <= 32'b00000111001110100110110000001100;
12'b011000000100: dataB <= 32'b00100000111111000000110111001010;
12'b011000000101: dataB <= 32'b00001010011000100001110101011100;
12'b011000000110: dataB <= 32'b00101100111110111010100100010000;
12'b011000000111: dataB <= 32'b00000111000100010000100010001100;
12'b011000001000: dataB <= 32'b11100111110001010011011010001011;
12'b011000001001: dataB <= 32'b00000010000110001100110101110110;
12'b011000001010: dataB <= 32'b01101000010101000000110101101010;
12'b011000001011: dataB <= 32'b00000110100001011010100101111001;
12'b011000001100: dataB <= 32'b11011000110100111010100111000111;
12'b011000001101: dataB <= 32'b00001001010111011011110111000000;
12'b011000001110: dataB <= 32'b01111101010010100011111100101101;
12'b011000001111: dataB <= 32'b00001110010111110001101011100101;
12'b011000010000: dataB <= 32'b10101101000100100001100011001101;
12'b011000010001: dataB <= 32'b00001100111011101001110010001100;
12'b011000010010: dataB <= 32'b01101010001011000011111111001111;
12'b011000010011: dataB <= 32'b00000110001100001110111101111000;
12'b011000010100: dataB <= 32'b11010101111011001011000011110110;
12'b011000010101: dataB <= 32'b00001010110010100001011101010110;
12'b011000010110: dataB <= 32'b10011110111101101010011001001000;
12'b011000010111: dataB <= 32'b00001010100010000100110110010010;
12'b011000011000: dataB <= 32'b11001001000111100100011100010100;
12'b011000011001: dataB <= 32'b00001101001000101110110000001011;
12'b011000011010: dataB <= 32'b00010001010000101010100000110000;
12'b011000011011: dataB <= 32'b00001001100001100010011101100100;
12'b011000011100: dataB <= 32'b11011111111001100000011001100010;
12'b011000011101: dataB <= 32'b00001011110101101101101111110011;
12'b011000011110: dataB <= 32'b00100100110001000011101011101000;
12'b011000011111: dataB <= 32'b00001000111101101101101110111010;
12'b011000100000: dataB <= 32'b11101011011100011001111010100101;
12'b011000100001: dataB <= 32'b00000001010111101010111111000100;
12'b011000100010: dataB <= 32'b10001111001010110011011001110001;
12'b011000100011: dataB <= 32'b00001110101110111101001110111001;
12'b011000100100: dataB <= 32'b01111011011101110110101100110101;
12'b011000100101: dataB <= 32'b00000101100001010010100010111101;
12'b011000100110: dataB <= 32'b00011101100100111000110110101001;
12'b011000100111: dataB <= 32'b00001001011110011001111010001101;
12'b011000101000: dataB <= 32'b01101000101100001010111001001101;
12'b011000101001: dataB <= 32'b00001110001011011111010001110011;
12'b011000101010: dataB <= 32'b10110000110000100001100101001000;
12'b011000101011: dataB <= 32'b00001000011011111101010001101100;
12'b011000101100: dataB <= 32'b11111000011100100011111100100101;
12'b011000101101: dataB <= 32'b00001001101001001111000101100011;
12'b011000101110: dataB <= 32'b10000101011010111100000100111101;
12'b011000101111: dataB <= 32'b00001000000111101010011010110010;
12'b011000110000: dataB <= 32'b11110011011101001010010010101101;
12'b011000110001: dataB <= 32'b00000100111001010111111010110100;
12'b011000110010: dataB <= 32'b10010001110110110001011001101001;
12'b011000110011: dataB <= 32'b00000011001110011110101101101110;
12'b011000110100: dataB <= 32'b11111010111011010100111111010001;
12'b011000110101: dataB <= 32'b00001011000010100110010110100100;
12'b011000110110: dataB <= 32'b01100000001110011011101000010010;
12'b011000110111: dataB <= 32'b00000111110111111001011110010000;
12'b011000111000: dataB <= 32'b01010011001111101011100100011100;
12'b011000111001: dataB <= 32'b00000100110010011101000100001101;
12'b011000111010: dataB <= 32'b11110001000010100100010101011000;
12'b011000111011: dataB <= 32'b00000110001000010000110111110010;
12'b011000111100: dataB <= 32'b00100101000001111001110110101100;
12'b011000111101: dataB <= 32'b00000000101011111000011111010010;
12'b011000111110: dataB <= 32'b01010000110001111100011110001100;
12'b011000111111: dataB <= 32'b00001001101000011110101110010000;
12'b011001000000: dataB <= 32'b10010101110010010101101011010100;
12'b011001000001: dataB <= 32'b00001110011000100001111011010100;
12'b011001000010: dataB <= 32'b10111000011110010001000111000111;
12'b011001000011: dataB <= 32'b00001001011010101101100001000100;
12'b011001000100: dataB <= 32'b00101110110100011101111110001011;
12'b011001000101: dataB <= 32'b00001101011010111011010101000101;
12'b011001000110: dataB <= 32'b01011001011010001100111111010001;
12'b011001000111: dataB <= 32'b00001011101110001011101011010011;
12'b011001001000: dataB <= 32'b01100010011100100001100000101011;
12'b011001001001: dataB <= 32'b00000100110011000111011101010000;
12'b011001001010: dataB <= 32'b01011111100111001100011010110101;
12'b011001001011: dataB <= 32'b00000110110101100111001111010100;
12'b011001001100: dataB <= 32'b10101000011101100001100000101111;
12'b011001001101: dataB <= 32'b00001101001000001101011010011000;
12'b011001001110: dataB <= 32'b10110100100010000001001010100011;
12'b011001001111: dataB <= 32'b00001000000001110000001110011010;
12'b011001010000: dataB <= 32'b01100001010010111000110000110100;
12'b011001010001: dataB <= 32'b00001011100010110010010110100100;
12'b011001010010: dataB <= 32'b00011000111010001101011011011101;
12'b011001010011: dataB <= 32'b00000110011101111011010010101010;
12'b011001010100: dataB <= 32'b11001100111010001000100010101010;
12'b011001010101: dataB <= 32'b00000111010111010101101011000000;
12'b011001010110: dataB <= 32'b11011000110110001110001010110110;
12'b011001010111: dataB <= 32'b00000010010010100110101100001010;
12'b011001011000: dataB <= 32'b11101110011101100101011000110010;
12'b011001011001: dataB <= 32'b00000111001110100100110000001100;
12'b011001011010: dataB <= 32'b01100000111110101000100110101010;
12'b011001011011: dataB <= 32'b00001011010110100111110001100100;
12'b011001011100: dataB <= 32'b00101010111010110010010100010001;
12'b011001011101: dataB <= 32'b00000110000101001110101010001100;
12'b011001011110: dataB <= 32'b11101101101101001011101001101010;
12'b011001011111: dataB <= 32'b00000001001001001100111110000110;
12'b011001100000: dataB <= 32'b10100010010000101001010101001011;
12'b011001100001: dataB <= 32'b00000101000001011000100101101001;
12'b011001100010: dataB <= 32'b10010110111000110011000110100111;
12'b011001100011: dataB <= 32'b00001001110111100001111010110000;
12'b011001100100: dataB <= 32'b11111101000110100011111100001011;
12'b011001100101: dataB <= 32'b00001111010101110101100011101100;
12'b011001100110: dataB <= 32'b10101100111100010010000011001111;
12'b011001100111: dataB <= 32'b00001101111001101101101110001100;
12'b011001101000: dataB <= 32'b01100100000111000011101110101100;
12'b011001101001: dataB <= 32'b00000110001100010001000101101000;
12'b011001101010: dataB <= 32'b00011011111011000010100100011000;
12'b011001101011: dataB <= 32'b00001010110001100101011101101111;
12'b011001101100: dataB <= 32'b01011110111101100010011000101000;
12'b011001101101: dataB <= 32'b00001001000001000011000010001010;
12'b011001101110: dataB <= 32'b10001001001111100011111100010011;
12'b011001101111: dataB <= 32'b00001100100110101100101000001100;
12'b011001110000: dataB <= 32'b01010011010100100011000000110010;
12'b011001110001: dataB <= 32'b00001000000001011110011101101100;
12'b011001110010: dataB <= 32'b01100101111001001000101000000010;
12'b011001110011: dataB <= 32'b00001100010011110001101011110011;
12'b011001110100: dataB <= 32'b11100010101101000011111010100111;
12'b011001110101: dataB <= 32'b00001010011101110001101010101001;
12'b011001110110: dataB <= 32'b01101101011000010010101001100101;
12'b011001110111: dataB <= 32'b00000010011001101010111011001100;
12'b011001111000: dataB <= 32'b01001111010010110011001001110001;
12'b011001111001: dataB <= 32'b00001110101011111101000010101001;
12'b011001111010: dataB <= 32'b11111101010010001110101101010011;
12'b011001111011: dataB <= 32'b00000100000010010000100111000100;
12'b011001111100: dataB <= 32'b00011111100100101001010110001001;
12'b011001111101: dataB <= 32'b00001010111110011111111010010101;
12'b011001111110: dataB <= 32'b01100110101000001011101000101101;
12'b011001111111: dataB <= 32'b00001101101001100001010001110011;
12'b011010000000: dataB <= 32'b10101110101100010010000100101001;
12'b011010000001: dataB <= 32'b00001001011010111101000101110100;
12'b011010000010: dataB <= 32'b00110100010100100100011011000011;
12'b011010000011: dataB <= 32'b00001001001001001111001001100100;
12'b011010000100: dataB <= 32'b01000111100010111011110110011110;
12'b011010000101: dataB <= 32'b00000111001000100110010110100010;
12'b011010000110: dataB <= 32'b10110101010100111010100010101111;
12'b011010000111: dataB <= 32'b00000101111010011011111010110100;
12'b011010001000: dataB <= 32'b10010111111010100001001001001001;
12'b011010001001: dataB <= 32'b00000011001111011110101101111110;
12'b011010001010: dataB <= 32'b10111010101111011100011111001110;
12'b011010001011: dataB <= 32'b00001010000001100010010010100100;
12'b011010001100: dataB <= 32'b01011010001110011011101000010010;
12'b011010001101: dataB <= 32'b00001000010111111101010101111000;
12'b011010001110: dataB <= 32'b11010101010011101010110101011110;
12'b011010001111: dataB <= 32'b00000100110011011111001000011101;
12'b011010010000: dataB <= 32'b00101110111010100100000110011001;
12'b011010010001: dataB <= 32'b00000101001001010000111011101010;
12'b011010010010: dataB <= 32'b10100101000001110001110110001101;
12'b011010010011: dataB <= 32'b00000000101110110100010111000001;
12'b011010010100: dataB <= 32'b01001110110101111100011101101010;
12'b011010010101: dataB <= 32'b00001001000111011110101101111000;
12'b011010010110: dataB <= 32'b00011001110110011101101011110010;
12'b011010010111: dataB <= 32'b00001110110101100111110111010100;
12'b011010011000: dataB <= 32'b11110100010110000000110110100111;
12'b011010011001: dataB <= 32'b00001010011001110001011101000100;
12'b011010011010: dataB <= 32'b01101100101100101110101101101001;
12'b011010011011: dataB <= 32'b00001110010111111101001001001101;
12'b011010011100: dataB <= 32'b11011011011010010100111111001110;
12'b011010011101: dataB <= 32'b00001011001101001111110011001010;
12'b011010011110: dataB <= 32'b11011110011100010010000000101110;
12'b011010011111: dataB <= 32'b00000101010100001011101001000000;
12'b011010100000: dataB <= 32'b10100011100111001011111010110100;
12'b011010100001: dataB <= 32'b00000111010110100111001111010011;
12'b011010100010: dataB <= 32'b10100110011101010001110000110010;
12'b011010100011: dataB <= 32'b00001100100110010001011110000000;
12'b011010100100: dataB <= 32'b01110000011001110001001001100010;
12'b011010100101: dataB <= 32'b00000110100001101010001010010010;
12'b011010100110: dataB <= 32'b00100001010010100000010001010111;
12'b011010100111: dataB <= 32'b00001010000001101100001110100100;
12'b011010101000: dataB <= 32'b11011000111010011101011100011100;
12'b011010101001: dataB <= 32'b00000111111101111101000110011001;
12'b011010101010: dataB <= 32'b10001101000001111000100010101100;
12'b011010101011: dataB <= 32'b00000111110111011001101110101000;
12'b011010101100: dataB <= 32'b10010110111010010110001011010100;
12'b011010101101: dataB <= 32'b00000010110100100100101100001011;
12'b011010101110: dataB <= 32'b10101010010101101101101000110010;
12'b011010101111: dataB <= 32'b00000110101111100010101100010101;
12'b011010110000: dataB <= 32'b01100000111110010000010110001011;
12'b011010110001: dataB <= 32'b00001011110101101011101101100100;
12'b011010110010: dataB <= 32'b00101010110010101001110100110010;
12'b011010110011: dataB <= 32'b00000101000110001100110010001100;
12'b011010110100: dataB <= 32'b10110001101001001100001001001001;
12'b011010110101: dataB <= 32'b00000000101100001101000110010110;
12'b011010110110: dataB <= 32'b11011110010000011001110100101100;
12'b011010110111: dataB <= 32'b00000100000011010110101001011001;
12'b011010111000: dataB <= 32'b01010110111100101011100101101000;
12'b011010111001: dataB <= 32'b00001010010110100101110110011000;
12'b011010111010: dataB <= 32'b00111100111010100011101011101001;
12'b011010111011: dataB <= 32'b00001111010010110111010111101100;
12'b011010111100: dataB <= 32'b01101100111000001010110011010000;
12'b011010111101: dataB <= 32'b00001110110111110001100110010100;
12'b011010111110: dataB <= 32'b10011110000111000011001110001001;
12'b011010111111: dataB <= 32'b00000101101101010001001001010000;
12'b011011000000: dataB <= 32'b00100001111010111010000101011001;
12'b011011000001: dataB <= 32'b00001010110000100111011001111111;
12'b011011000010: dataB <= 32'b01011110111101011010100111101000;
12'b011011000011: dataB <= 32'b00000111100001000101001010000010;
12'b011011000100: dataB <= 32'b01001011010111011011001100110001;
12'b011011000101: dataB <= 32'b00001011100101101010100100001101;
12'b011011000110: dataB <= 32'b01010101011000011011110001010101;
12'b011011000111: dataB <= 32'b00000110100001011010011101101100;
12'b011011001000: dataB <= 32'b10101001111000111000110110100010;
12'b011011001001: dataB <= 32'b00001100010001110101100011101010;
12'b011011001010: dataB <= 32'b10100000101101000100011010000110;
12'b011011001011: dataB <= 32'b00001011011100110101100010100001;
12'b011011001100: dataB <= 32'b11101111010000001011011000100100;
12'b011011001101: dataB <= 32'b00000011011011101000110111001011;
12'b011011001110: dataB <= 32'b00010001010110101010111001110000;
12'b011011001111: dataB <= 32'b00001110001001111100110110011001;
12'b011011010000: dataB <= 32'b01111101000110011110101101010001;
12'b011011010001: dataB <= 32'b00000011000100001110101111000100;
12'b011011010010: dataB <= 32'b11100011100100011010000101101010;
12'b011011010011: dataB <= 32'b00001011111100100101111010011100;
12'b011011010100: dataB <= 32'b10100100101000001100011000101101;
12'b011011010101: dataB <= 32'b00001100100111100011010001101011;
12'b011011010110: dataB <= 32'b10101100100100001010110100001011;
12'b011011010111: dataB <= 32'b00001010011010111100111001110100;
12'b011011011000: dataB <= 32'b01101110001100101100111010000010;
12'b011011011001: dataB <= 32'b00001000001000010001010001100100;
12'b011011011010: dataB <= 32'b00001011101010110011010111111110;
12'b011011011011: dataB <= 32'b00000110101000100010010110011010;
12'b011011011100: dataB <= 32'b00110111001100111011000010110001;
12'b011011011101: dataB <= 32'b00000110111010100001111010111100;
12'b011011011110: dataB <= 32'b10011101111010010000111000001000;
12'b011011011111: dataB <= 32'b00000011010001011100101110001110;
12'b011011100000: dataB <= 32'b01111000100111011011101111001011;
12'b011011100001: dataB <= 32'b00001000100001011100010010101100;
12'b011011100010: dataB <= 32'b01010110010010011011011000010010;
12'b011011100011: dataB <= 32'b00001001010110111101001001100000;
12'b011011100100: dataB <= 32'b10010111010111100010010110111110;
12'b011011100101: dataB <= 32'b00000101010100011111001000101110;
12'b011011100110: dataB <= 32'b10101110110110100011110111011010;
12'b011011100111: dataB <= 32'b00000100101010010001000011011001;
12'b011011101000: dataB <= 32'b00100100111101100001110110001110;
12'b011011101001: dataB <= 32'b00000000110001101110001110110001;
12'b011011101010: dataB <= 32'b01001110111110000100011101000111;
12'b011011101011: dataB <= 32'b00001000000111011100101101100000;
12'b011011101100: dataB <= 32'b10011111110110100101011011110001;
12'b011011101101: dataB <= 32'b00001111010010101101110011010011;
12'b011011101110: dataB <= 32'b00101110001101110001000101101000;
12'b011011101111: dataB <= 32'b00001010111000110011010101001101;
12'b011011110000: dataB <= 32'b10101010101000111111001100100111;
12'b011011110001: dataB <= 32'b00001111010101111100111101010101;
12'b011011110010: dataB <= 32'b10011111011110011100101111001011;
12'b011011110011: dataB <= 32'b00001010101011010011110111000010;
12'b011011110100: dataB <= 32'b01011010011100001010110000110001;
12'b011011110101: dataB <= 32'b00000101110101001111110000101001;
12'b011011110110: dataB <= 32'b00100111100011001011011011010010;
12'b011011110111: dataB <= 32'b00000111110110101001001011010011;
12'b011011111000: dataB <= 32'b10100010011001000010000000110101;
12'b011011111001: dataB <= 32'b00001011100101010011100101101000;
12'b011011111010: dataB <= 32'b01101100010001100001011000000010;
12'b011011111011: dataB <= 32'b00000101000001100100000110001010;
12'b011011111100: dataB <= 32'b11100011010010010000010010011001;
12'b011011111101: dataB <= 32'b00001000100001101000001010100011;
12'b011011111110: dataB <= 32'b11011000111110100101001101011010;
12'b011011111111: dataB <= 32'b00001001011101111100111010001001;
12'b011100000000: dataB <= 32'b01001101001001100000100010001110;
12'b011100000001: dataB <= 32'b00001000110111011111110010010000;
12'b011100000010: dataB <= 32'b01010110111110100101111011110011;
12'b011100000011: dataB <= 32'b00000011010110100010101000001100;
12'b011100000100: dataB <= 32'b00100110010001110101101001010001;
12'b011100000101: dataB <= 32'b00000110101111100000101100011110;
12'b011100000110: dataB <= 32'b10100000111101111000010101101100;
12'b011100000111: dataB <= 32'b00001100010100110001101001100100;
12'b011100001000: dataB <= 32'b11101000101110011001110101010100;
12'b011100001001: dataB <= 32'b00000100000111001010111010001011;
12'b011100001010: dataB <= 32'b10110101100001001100011000101001;
12'b011100001011: dataB <= 32'b00000000101111001111001110100110;
12'b011100001100: dataB <= 32'b00011010010000010010010100001101;
12'b011100001101: dataB <= 32'b00000010100101010100101101001010;
12'b011100001110: dataB <= 32'b01010110111100101100000101001001;
12'b011100001111: dataB <= 32'b00001011010101101011110110000000;
12'b011100010000: dataB <= 32'b10111100101110011011011011001000;
12'b011100010001: dataB <= 32'b00001111001111111001001111101011;
12'b011100010010: dataB <= 32'b01101010110100001011100011010010;
12'b011100010011: dataB <= 32'b00001111010100110101011110010100;
12'b011100010100: dataB <= 32'b11011000000110111010101101100111;
12'b011100010101: dataB <= 32'b00000101101110010011010000111000;
12'b011100010110: dataB <= 32'b00100111111010101001110110011010;
12'b011100010111: dataB <= 32'b00001010101111101001010110010111;
12'b011100011000: dataB <= 32'b01011110111101010010110111001000;
12'b011100011001: dataB <= 32'b00000110000001000101010101110010;
12'b011100011010: dataB <= 32'b11001111011111010010101100101111;
12'b011100011011: dataB <= 32'b00001010100100100110100000011101;
12'b011100011100: dataB <= 32'b10010111011100011100010001111000;
12'b011100011101: dataB <= 32'b00000101100001011000100001101100;
12'b011100011110: dataB <= 32'b11101111110000101001010101100011;
12'b011100011111: dataB <= 32'b00001100010000110111011011100001;
12'b011100100000: dataB <= 32'b01100000101101000100101001000101;
12'b011100100001: dataB <= 32'b00001100111010110111011010010001;
12'b011100100010: dataB <= 32'b10110001001100001011110111100100;
12'b011100100011: dataB <= 32'b00000100011101101000110011001011;
12'b011100100100: dataB <= 32'b11010011011010100010101001101111;
12'b011100100101: dataB <= 32'b00001101000110111010101010000000;
12'b011100100110: dataB <= 32'b00111100111010101110011101001110;
12'b011100100111: dataB <= 32'b00000010000110001100110111000100;
12'b011100101000: dataB <= 32'b11100111100000001010100101001011;
12'b011100101001: dataB <= 32'b00001101011010101011110110011100;
12'b011100101010: dataB <= 32'b10100010100100001101001000001100;
12'b011100101011: dataB <= 32'b00001011100101100101010001101011;
12'b011100101100: dataB <= 32'b11101010100000001011100011101100;
12'b011100101101: dataB <= 32'b00001011011001111100101101111100;
12'b011100101110: dataB <= 32'b01101010000100101101011000100010;
12'b011100101111: dataB <= 32'b00000111101000010011010101100100;
12'b011100110000: dataB <= 32'b00010001110010110011001001011110;
12'b011100110001: dataB <= 32'b00000101101001011100010110010010;
12'b011100110010: dataB <= 32'b11111001000000110011100011010011;
12'b011100110011: dataB <= 32'b00000111111011100111111010111011;
12'b011100110100: dataB <= 32'b01100011111001111000110111101000;
12'b011100110101: dataB <= 32'b00000011110011011010110010011110;
12'b011100110110: dataB <= 32'b00110100011011010011001110101001;
12'b011100110111: dataB <= 32'b00000111000001011000010110101100;
12'b011100111000: dataB <= 32'b10010010010110010011001000110001;
12'b011100111001: dataB <= 32'b00001001110110111100111101001000;
12'b011100111010: dataB <= 32'b00011001011011010001101000011110;
12'b011100111011: dataB <= 32'b00000101110101011111001000111111;
12'b011100111100: dataB <= 32'b00101100101110100011101000011010;
12'b011100111101: dataB <= 32'b00000100001100010001000111001001;
12'b011100111110: dataB <= 32'b11100100111101010010000110001110;
12'b011100111111: dataB <= 32'b00000000110100101010000110100000;
12'b011101000000: dataB <= 32'b10001111000110000100011100000101;
12'b011101000001: dataB <= 32'b00000111000111011010110001001000;
12'b011101000010: dataB <= 32'b00100011110110101101001100001111;
12'b011101000011: dataB <= 32'b00001111010000110001101111001011;
12'b011101000100: dataB <= 32'b10101010000101011001000101001001;
12'b011101000101: dataB <= 32'b00001011110111110101001101010101;
12'b011101000110: dataB <= 32'b11101000100101001111011011100101;
12'b011101000111: dataB <= 32'b00001111010010111100110001011101;
12'b011101001000: dataB <= 32'b00100001011110011100011110101001;
12'b011101001001: dataB <= 32'b00001010101010011001111010111010;
12'b011101001010: dataB <= 32'b11011000100000001011100000110100;
12'b011101001011: dataB <= 32'b00000110010110010011110100011001;
12'b011101001100: dataB <= 32'b10101001100011001010111011110001;
12'b011101001101: dataB <= 32'b00001000110110101001000111001010;
12'b011101001110: dataB <= 32'b11011110011000111010100001110111;
12'b011101001111: dataB <= 32'b00001010100100010111101001011000;
12'b011101010000: dataB <= 32'b01101000001101010001010111000010;
12'b011101010001: dataB <= 32'b00000100000011011110000110000010;
12'b011101010010: dataB <= 32'b10100101001101111000010011011011;
12'b011101010011: dataB <= 32'b00000111000001100010001010100011;
12'b011101010100: dataB <= 32'b11011001000010100100111110010111;
12'b011101010101: dataB <= 32'b00001010011100111010101110000001;
12'b011101010110: dataB <= 32'b01001101010001010000110010010000;
12'b011101010111: dataB <= 32'b00001001010111100011110010000000;
12'b011101011000: dataB <= 32'b00010110111110101101101011110010;
12'b011101011001: dataB <= 32'b00000100011000100000101000001101;
12'b011101011010: dataB <= 32'b10100010010001111101101001010001;
12'b011101011011: dataB <= 32'b00000110101111100000101100101110;
12'b011101011100: dataB <= 32'b11100000111101100000010101001101;
12'b011101011101: dataB <= 32'b00001100010010110101100001101100;
12'b011101011110: dataB <= 32'b11100110101110001001100101010101;
12'b011101011111: dataB <= 32'b00000011101001001011000010001011;
12'b011101100000: dataB <= 32'b01110111011001010100101000001001;
12'b011101100001: dataB <= 32'b00000000110010001111010010110110;
12'b011101100010: dataB <= 32'b01010110010100001011000100001111;
12'b011101100011: dataB <= 32'b00000001100111010010110001000010;
12'b011101100100: dataB <= 32'b01010111000000101100100100101010;
12'b011101100101: dataB <= 32'b00001011110100101111101101101000;
12'b011101100110: dataB <= 32'b11111010100010011011001010000111;
12'b011101100111: dataB <= 32'b00001111001100111011000011100010;
12'b011101101000: dataB <= 32'b00101010110000001100010011110100;
12'b011101101001: dataB <= 32'b00001111010001110111010110010100;
12'b011101101010: dataB <= 32'b01010100001010110010011100100101;
12'b011101101011: dataB <= 32'b00000101001111010101010100101001;
12'b011101101100: dataB <= 32'b11101101110110011001100111011011;
12'b011101101101: dataB <= 32'b00001010101110101011010010100110;
12'b011101101110: dataB <= 32'b10011110111101001011010110001000;
12'b011101101111: dataB <= 32'b00000101000010001001011101101010;
12'b011101110000: dataB <= 32'b10010001100111001010001100101101;
12'b011101110001: dataB <= 32'b00001001000011100100100000100110;
12'b011101110010: dataB <= 32'b10011011100000100100110010111010;
12'b011101110011: dataB <= 32'b00000100000011010100100101110100;
12'b011101110100: dataB <= 32'b01110011101100011010000100100100;
12'b011101110101: dataB <= 32'b00001100001110111001001111010001;
12'b011101110110: dataB <= 32'b01011110101101001101001000000101;
12'b011101110111: dataB <= 32'b00001101011000111001001110000001;
12'b011101111000: dataB <= 32'b00110001000100001100100110100100;
12'b011101111001: dataB <= 32'b00000101111110100110101111000011;
12'b011101111010: dataB <= 32'b00010111100010010010011001101110;
12'b011101111011: dataB <= 32'b00001100000101111000011101110001;
12'b011101111100: dataB <= 32'b10111100101110110110001101001100;
12'b011101111101: dataB <= 32'b00000001001000001010111111000011;
12'b011101111110: dataB <= 32'b10101001011100001011010100101101;
12'b011101111111: dataB <= 32'b00001110011000110001110010100100;
12'b011110000000: dataB <= 32'b11011110100100010101110111101100;
12'b011110000001: dataB <= 32'b00001010100100100101010001101011;
12'b011110000010: dataB <= 32'b11100110011100001100010011101110;
12'b011110000011: dataB <= 32'b00001100010111111010100010000100;
12'b011110000100: dataB <= 32'b10100100000100111101110111000010;
12'b011110000101: dataB <= 32'b00000110101001010101011001101100;
12'b011110000110: dataB <= 32'b11010101111010101010111010011110;
12'b011110000111: dataB <= 32'b00000101001010011000010110000001;
12'b011110001000: dataB <= 32'b01110110111000110100000011010101;
12'b011110001001: dataB <= 32'b00001000111011101101110110110011;
12'b011110001010: dataB <= 32'b01101001111001101000110110101001;
12'b011110001011: dataB <= 32'b00000100010100011000110010101110;
12'b011110001100: dataB <= 32'b11110000010111001010101101100110;
12'b011110001101: dataB <= 32'b00000101100001010100011010101011;
12'b011110001110: dataB <= 32'b00001110011110010011001000110001;
12'b011110001111: dataB <= 32'b00001010010101111100110000110001;
12'b011110010000: dataB <= 32'b01011011011011000001011001111110;
12'b011110010001: dataB <= 32'b00000110110110100001001001001111;
12'b011110010010: dataB <= 32'b10101010101010011011101001011010;
12'b011110010011: dataB <= 32'b00000100001101010001001110111000;
12'b011110010100: dataB <= 32'b10100100111001001010010101101111;
12'b011110010101: dataB <= 32'b00000001010111100100000110001000;
12'b011110010110: dataB <= 32'b00001111001010000100011011000100;
12'b011110010111: dataB <= 32'b00000110100111011000110000110001;
12'b011110011000: dataB <= 32'b10101001110010110100101011101110;
12'b011110011001: dataB <= 32'b00001111001101110101100111001010;
12'b011110011010: dataB <= 32'b11100100000101001001010100101010;
12'b011110011011: dataB <= 32'b00001100010101110111000101011101;
12'b011110011100: dataB <= 32'b00100110100001100111101010100100;
12'b011110011101: dataB <= 32'b00001111001111111010101001101110;
12'b011110011110: dataB <= 32'b11100101011010011100011101100110;
12'b011110011111: dataB <= 32'b00001001101001011111111010101001;
12'b011110100000: dataB <= 32'b01010100100100001100010001010111;
12'b011110100001: dataB <= 32'b00000110110110011001111000010010;
12'b011110100010: dataB <= 32'b01101101011111000010101011110000;
12'b011110100011: dataB <= 32'b00001001010101101011000011000010;
12'b011110100100: dataB <= 32'b00011010011000110011000010011010;
12'b011110100101: dataB <= 32'b00001001000011011011101001001001;
12'b011110100110: dataB <= 32'b01100010001001000001110101100011;
12'b011110100111: dataB <= 32'b00000010100100011010000101110010;
12'b011110101000: dataB <= 32'b10100111001101100000010100011101;
12'b011110101001: dataB <= 32'b00000101100001011100001010011011;
12'b011110101010: dataB <= 32'b11011001000110101100101111010101;
12'b011110101011: dataB <= 32'b00001011011011111000100101110001;
12'b011110101100: dataB <= 32'b01001111010100111001010010010010;
12'b011110101101: dataB <= 32'b00001010010110100111101101101000;
12'b011110101110: dataB <= 32'b11010111000010110101011100010000;
12'b011110101111: dataB <= 32'b00000100111001011110101000010101;
12'b011110110000: dataB <= 32'b00011110010010001101101001010000;
12'b011110110001: dataB <= 32'b00000110110000011110101101000111;
12'b011110110010: dataB <= 32'b11100000111101010000100101001110;
12'b011110110011: dataB <= 32'b00001100110000110111011001101100;
12'b011110110100: dataB <= 32'b11100100101001111001100110010110;
12'b011110110101: dataB <= 32'b00000011001010001011001010001011;
12'b011110110110: dataB <= 32'b11111001001101010100110111001001;
12'b011110110111: dataB <= 32'b00000000110100010001011011000101;
12'b011110111000: dataB <= 32'b11010010011000001011110100010000;
12'b011110111001: dataB <= 32'b00000001001001010010110100111010;
12'b011110111010: dataB <= 32'b01010111000100110101000100001100;
12'b011110111011: dataB <= 32'b00001011110010110101101001011000;
12'b011110111100: dataB <= 32'b01110110011010010011001001000110;
12'b011110111101: dataB <= 32'b00001110101001111010111011011010;
12'b011110111110: dataB <= 32'b00101000101100001101000100010110;
12'b011110111111: dataB <= 32'b00001111001110111001001110010100;
12'b011111000000: dataB <= 32'b11001110001110100010001011100011;
12'b011111000001: dataB <= 32'b00000101010000010111011000011001;
12'b011111000010: dataB <= 32'b10110001110010001001101000011011;
12'b011111000011: dataB <= 32'b00001010101101101101001110110110;
12'b011111000100: dataB <= 32'b10011110111101001011100101101001;
12'b011111000101: dataB <= 32'b00000011100011001011101001100010;
12'b011111000110: dataB <= 32'b00010101101010111001101100001011;
12'b011111000111: dataB <= 32'b00001000000010100000100000111111;
12'b011111001000: dataB <= 32'b10011111100000101101010011111100;
12'b011111001001: dataB <= 32'b00000011000100010010101001110100;
12'b011111001010: dataB <= 32'b11110111100100001010100011000110;
12'b011111001011: dataB <= 32'b00001100001100111001000111000000;
12'b011111001100: dataB <= 32'b01011100101101010101010110100101;
12'b011111001101: dataB <= 32'b00001110010110111001000101101001;
12'b011111001110: dataB <= 32'b10110010111100010101010101100101;
12'b011111001111: dataB <= 32'b00000111011110100100101110111010;
12'b011111010000: dataB <= 32'b00011011100010001010011001101110;
12'b011111010001: dataB <= 32'b00001011000011110100010101100001;
12'b011111010010: dataB <= 32'b00111010100011000101101100101010;
12'b011111010011: dataB <= 32'b00000000101011001011000111000011;
12'b011111010100: dataB <= 32'b01101101011000001100000100101110;
12'b011111010101: dataB <= 32'b00001110110110110101101010100100;
12'b011111010110: dataB <= 32'b11011100100100100110010111101100;
12'b011111010111: dataB <= 32'b00001001100011100111001101101011;
12'b011111011000: dataB <= 32'b11100010011100001101000011010000;
12'b011111011001: dataB <= 32'b00001100110101110110011010000100;
12'b011111011010: dataB <= 32'b10011110000101001110010110000010;
12'b011111011011: dataB <= 32'b00000110001001011001011101101100;
12'b011111011100: dataB <= 32'b11011011111010100010101011111100;
12'b011111011101: dataB <= 32'b00000100101011010100011001110001;
12'b011111011110: dataB <= 32'b00110110110000110100100100010111;
12'b011111011111: dataB <= 32'b00001001111010110001101110110011;
12'b011111100000: dataB <= 32'b11101111110101011001000110001001;
12'b011111100001: dataB <= 32'b00000100110110011000110110111101;
12'b011111100010: dataB <= 32'b10101100001111000010001100100100;
12'b011111100011: dataB <= 32'b00000100000010010000011110101011;
12'b011111100100: dataB <= 32'b01001010100010001011001000110001;
12'b011111100101: dataB <= 32'b00001010110100111010100100100001;
12'b011111100110: dataB <= 32'b10011111011010110000111011011101;
12'b011111100111: dataB <= 32'b00000111010110100001001001100111;
12'b011111101000: dataB <= 32'b01101000100110011011011010011001;
12'b011111101001: dataB <= 32'b00000100001111010011010010100000;
12'b011111101010: dataB <= 32'b10100100111001000010110101110000;
12'b011111101011: dataB <= 32'b00000010011001011110000101111000;
12'b011111101100: dataB <= 32'b01010001010010000100011010000011;
12'b011111101101: dataB <= 32'b00000101101000011000110100100001;
12'b011111101110: dataB <= 32'b00101101101110110100011011101100;
12'b011111101111: dataB <= 32'b00001110101010111001011110111010;
12'b011111110000: dataB <= 32'b11011110000100111001110100001100;
12'b011111110001: dataB <= 32'b00001100110011110110111101101101;
12'b011111110010: dataB <= 32'b00100010100001111111101001100011;
12'b011111110011: dataB <= 32'b00001111001100111000011101111110;
12'b011111110100: dataB <= 32'b10100111011010011100001100100100;
12'b011111110101: dataB <= 32'b00001001001001100101111010011001;
12'b011111110110: dataB <= 32'b00010010101000001101000010011001;
12'b011111110111: dataB <= 32'b00000111110110011111111000001011;
12'b011111111000: dataB <= 32'b11101111010110110010001011101110;
12'b011111111001: dataB <= 32'b00001001110101101010111110110001;
12'b011111111010: dataB <= 32'b10010110011100110011100011111100;
12'b011111111011: dataB <= 32'b00001000000010011111101100110001;
12'b011111111100: dataB <= 32'b01011110001000110010010100100100;
12'b011111111101: dataB <= 32'b00000001100111010100001001101010;
12'b011111111110: dataB <= 32'b01100111001001001000100101111110;
12'b011111111111: dataB <= 32'b00000100000010011000001010011011;
12'b100000000000: dataB <= 32'b11011001000110101100011111010010;
12'b100000000001: dataB <= 32'b00001100111001110100011101100001;
12'b100000000010: dataB <= 32'b10010011011100101001100010110100;
12'b100000000011: dataB <= 32'b00001010110101101011101001010000;
12'b100000000100: dataB <= 32'b01010111000110111100111100001110;
12'b100000000101: dataB <= 32'b00000101111010011100101000100110;
12'b100000000110: dataB <= 32'b10011010010010010101101001010000;
12'b100000000111: dataB <= 32'b00000110110000011100101101010111;
12'b100000001000: dataB <= 32'b11100000111100111000110101001111;
12'b100000001001: dataB <= 32'b00001100101110111001010001110100;
12'b100000001010: dataB <= 32'b11100010101001101001100110110110;
12'b100000001011: dataB <= 32'b00000010101100001101010010001011;
12'b100000001100: dataB <= 32'b01111001000101011101000110101001;
12'b100000001101: dataB <= 32'b00000001110111010101011111001101;
12'b100000001110: dataB <= 32'b01001110100000001100100100010010;
12'b100000001111: dataB <= 32'b00000000101100010010111100110011;
12'b100000010000: dataB <= 32'b00100011010010100110010110010111;
12'b100000010001: dataB <= 32'b00001001001000110100010100001101;
12'b100000010010: dataB <= 32'b00001100010001100011010011001101;
12'b100000010011: dataB <= 32'b00000100100010011100001001001001;
12'b100000010100: dataB <= 32'b01010110101110100111101011010111;
12'b100000010101: dataB <= 32'b00000111000001100110001110000011;
12'b100000010110: dataB <= 32'b00000111100001000010110001101000;
12'b100000010111: dataB <= 32'b00001000010101101101010000111111;
12'b100000011000: dataB <= 32'b01111000011100110011101101101111;
12'b100000011001: dataB <= 32'b00000110101010100110100111010010;
12'b100000011010: dataB <= 32'b11011111000001110101100100110100;
12'b100000011011: dataB <= 32'b00000001111000110101101001010100;
12'b100000011100: dataB <= 32'b00110101010100110010000101100111;
12'b100000011101: dataB <= 32'b00000001001111010000111111100110;
12'b100000011110: dataB <= 32'b01110001000010101110101110011000;
12'b100000011111: dataB <= 32'b00000010011001010101011010010100;
12'b100000100000: dataB <= 32'b11110010010001010111100011011001;
12'b100000100001: dataB <= 32'b00000110000111100010001100011001;
12'b100000100010: dataB <= 32'b10010111000110101101010010110010;
12'b100000100011: dataB <= 32'b00001011000011100010001100101100;
12'b100000100100: dataB <= 32'b00011110011010101111010010110100;
12'b100000100101: dataB <= 32'b00001111010001010110110101010010;
12'b100000100110: dataB <= 32'b11110001001001001011100111001100;
12'b100000100111: dataB <= 32'b00000001101001001010010100100100;
12'b100000101000: dataB <= 32'b11010000001010110001110101000110;
12'b100000101001: dataB <= 32'b00000101111110100011101001100001;
12'b100000101010: dataB <= 32'b11101100100110000111100111010110;
12'b100000101011: dataB <= 32'b00001011000010110100010110001010;
12'b100000101100: dataB <= 32'b10010011000111001110110110010000;
12'b100000101101: dataB <= 32'b00000001101100100110110001111100;
12'b100000101110: dataB <= 32'b11001110111010100111101000011001;
12'b100000101111: dataB <= 32'b00001010100110001100010010011011;
12'b100000110000: dataB <= 32'b10000011000011001101100001010011;
12'b100000110001: dataB <= 32'b00000100110011101111001110010100;
12'b100000110010: dataB <= 32'b01111101001001010010111110001000;
12'b100000110011: dataB <= 32'b00000101110110001101010100111100;
12'b100000110100: dataB <= 32'b01011000010010010110011011110111;
12'b100000110101: dataB <= 32'b00001101001100110110011101100010;
12'b100000110110: dataB <= 32'b00111010100000100101000100110011;
12'b100000110111: dataB <= 32'b00001011010110011011001110111010;
12'b100000111000: dataB <= 32'b10000110100101000001110010000110;
12'b100000111001: dataB <= 32'b00000001010111001111011101110010;
12'b100000111010: dataB <= 32'b11010001101001100011101000101110;
12'b100000111011: dataB <= 32'b00001010001010010010001000101110;
12'b100000111100: dataB <= 32'b11101101000000011010011110101001;
12'b100000111101: dataB <= 32'b00001011010001100100111111110100;
12'b100000111110: dataB <= 32'b11010010101101101011001100101011;
12'b100000111111: dataB <= 32'b00000111110111101001011000001010;
12'b100001000000: dataB <= 32'b00011100110101011101111000010100;
12'b100001000001: dataB <= 32'b00001100111011000011000000010100;
12'b100001000010: dataB <= 32'b11101001011110001011110001101011;
12'b100001000011: dataB <= 32'b00000100010100011011001100101110;
12'b100001000100: dataB <= 32'b00110110100110001010010110001000;
12'b100001000101: dataB <= 32'b00000101000010101110001101000010;
12'b100001000110: dataB <= 32'b10000011000000111110000110010111;
12'b100001000111: dataB <= 32'b00001001100110011110010010111100;
12'b100001001000: dataB <= 32'b00010000111011110100000001101100;
12'b100001001001: dataB <= 32'b00000110000001001110001111000100;
12'b100001001010: dataB <= 32'b00101100110010000011000010000110;
12'b100001001011: dataB <= 32'b00000100101101111100110100110011;
12'b100001001100: dataB <= 32'b10010101011010100111101100111011;
12'b100001001101: dataB <= 32'b00001011010000111101000001100111;
12'b100001001110: dataB <= 32'b01101010100001000010010111001000;
12'b100001001111: dataB <= 32'b00001010101100011110101000111010;
12'b100001010000: dataB <= 32'b01001111010001110110011110011000;
12'b100001010001: dataB <= 32'b00000001001111110111000000110110;
12'b100001010010: dataB <= 32'b10000101000001001110010010010110;
12'b100001010011: dataB <= 32'b00000011111100000101010101001100;
12'b100001010100: dataB <= 32'b00100100110000010101101111010100;
12'b100001010101: dataB <= 32'b00000001010111000101001101101011;
12'b100001010110: dataB <= 32'b11100011001110001010101001000001;
12'b100001010111: dataB <= 32'b00001100100110001110010100111100;
12'b100001011000: dataB <= 32'b01101111011000110110101010011010;
12'b100001011001: dataB <= 32'b00001010101010110100101000010101;
12'b100001011010: dataB <= 32'b11100011010010011010000111000111;
12'b100001011011: dataB <= 32'b00001101010100010101000111001110;
12'b100001011100: dataB <= 32'b01001001001010110011011000001101;
12'b100001011101: dataB <= 32'b00001000010010010111000111110101;
12'b100001011110: dataB <= 32'b01011110111100011110000111110101;
12'b100001011111: dataB <= 32'b00000111000110101000001110011100;
12'b100001100000: dataB <= 32'b10010100111000110100101011010010;
12'b100001100001: dataB <= 32'b00000110011010101001100101111011;
12'b100001100010: dataB <= 32'b10100010001110100101000100110010;
12'b100001100011: dataB <= 32'b00001011111100101111010110101001;
12'b100001100100: dataB <= 32'b01010001100010010111101001010111;
12'b100001100101: dataB <= 32'b00000110011110011111011001101110;
12'b100001100110: dataB <= 32'b10100001010010010110100101010110;
12'b100001100111: dataB <= 32'b00001010001000110110100000001100;
12'b100001101000: dataB <= 32'b11010000001001100011000011101011;
12'b100001101001: dataB <= 32'b00000110000001100000001001011000;
12'b100001101010: dataB <= 32'b01011000101010001111101010011000;
12'b100001101011: dataB <= 32'b00001000100001101010010010000011;
12'b100001101100: dataB <= 32'b10000101010101001010010010100110;
12'b100001101101: dataB <= 32'b00000111110101101011010100101110;
12'b100001101110: dataB <= 32'b11111010100100110011001101110001;
12'b100001101111: dataB <= 32'b00000111001010101000101011011010;
12'b100001110000: dataB <= 32'b10011111000001101101100100010011;
12'b100001110001: dataB <= 32'b00000001010101101111101101010100;
12'b100001110010: dataB <= 32'b11110011011101000001100110100110;
12'b100001110011: dataB <= 32'b00000001101101010000110111010110;
12'b100001110100: dataB <= 32'b01110001001010011110111101011010;
12'b100001110101: dataB <= 32'b00000001110111010011010110010100;
12'b100001110110: dataB <= 32'b01110110011001000111000010010110;
12'b100001110111: dataB <= 32'b00000111000111100110001100101001;
12'b100001111000: dataB <= 32'b11010111000010100101100010101111;
12'b100001111001: dataB <= 32'b00001100000101100110001100101011;
12'b100001111010: dataB <= 32'b11100010011110010111100010010010;
12'b100001111011: dataB <= 32'b00001111010100010110110001100001;
12'b100001111100: dataB <= 32'b01110001010001001011010111001100;
12'b100001111101: dataB <= 32'b00000010100111001110001100100100;
12'b100001111110: dataB <= 32'b11010110000111000010010110000101;
12'b100001111111: dataB <= 32'b00000100011101011111101001110001;
12'b100010000000: dataB <= 32'b11101110101101101111100110110110;
12'b100010000001: dataB <= 32'b00001100000011111000011110010010;
12'b100010000010: dataB <= 32'b10010011000010111111010110010000;
12'b100010000011: dataB <= 32'b00000010001010101000110101111100;
12'b100010000100: dataB <= 32'b11001110110010001111100111011000;
12'b100010000101: dataB <= 32'b00001011100111010000001010011011;
12'b100010000110: dataB <= 32'b10000010110110111110000001010001;
12'b100010000111: dataB <= 32'b00000100110010101101010110010100;
12'b100010001000: dataB <= 32'b11111101010101011010101111001011;
12'b100010001001: dataB <= 32'b00000101010101001011001100111011;
12'b100010001010: dataB <= 32'b01011100010010000110011010111001;
12'b100010001011: dataB <= 32'b00001101101110111010100101101010;
12'b100010001100: dataB <= 32'b10111100101100011100100100110010;
12'b100010001101: dataB <= 32'b00001010010111011001001111001010;
12'b100010001110: dataB <= 32'b10001010011101010001100011000100;
12'b100010001111: dataB <= 32'b00000000110100001101010101111010;
12'b100010010000: dataB <= 32'b01001111100001100011011000101110;
12'b100010010001: dataB <= 32'b00001010101011011000000100100110;
12'b100010010010: dataB <= 32'b10101101001000101001111111001100;
12'b100010010011: dataB <= 32'b00001011010010100100111111101101;
12'b100010010100: dataB <= 32'b00010100101001110011001101001101;
12'b100010010101: dataB <= 32'b00000110110111100111011100010010;
12'b100010010110: dataB <= 32'b10011100110101001101100111110100;
12'b100010010111: dataB <= 32'b00001011111101000010110100010011;
12'b100010011000: dataB <= 32'b01100101100010001011110010001001;
12'b100010011001: dataB <= 32'b00000011110010011001001100100110;
12'b100010011010: dataB <= 32'b10111000101110010010010111001000;
12'b100010011011: dataB <= 32'b00000110100001110010010101010001;
12'b100010011100: dataB <= 32'b00000010110100101101100101010110;
12'b100010011101: dataB <= 32'b00001010100111100010010010111101;
12'b100010011110: dataB <= 32'b10010000110011110100110010001010;
12'b100010011111: dataB <= 32'b00000111100001010100001011000100;
12'b100010100000: dataB <= 32'b10101100110110001011000011000100;
12'b100010100001: dataB <= 32'b00000100101100111101000000111010;
12'b100010100010: dataB <= 32'b01010011010110001111101011111101;
12'b100010100011: dataB <= 32'b00001011010010111101001101001111;
12'b100010100100: dataB <= 32'b11101110100101010001111000001000;
12'b100010100101: dataB <= 32'b00001010101101100000101001001001;
12'b100010100110: dataB <= 32'b10001101001001100110011101011011;
12'b100010100111: dataB <= 32'b00000001101101110101001000100101;
12'b100010101000: dataB <= 32'b01000100111000111101110001110100;
12'b100010101001: dataB <= 32'b00000010011010000011001001001100;
12'b100010101010: dataB <= 32'b00100110110000001100111110110111;
12'b100010101011: dataB <= 32'b00000000110100000101000101110011;
12'b100010101100: dataB <= 32'b01100011001110010010101010100001;
12'b100010101101: dataB <= 32'b00001101101001010010001100111100;
12'b100010101110: dataB <= 32'b10101011100000101110001001011011;
12'b100010101111: dataB <= 32'b00001011001011110110110000001100;
12'b100010110000: dataB <= 32'b01100001010010101010011000000111;
12'b100010110001: dataB <= 32'b00001100110110010101000010111111;
12'b100010110010: dataB <= 32'b11001001000010110011101000001101;
12'b100010110011: dataB <= 32'b00001000010010010111000011100101;
12'b100010110100: dataB <= 32'b10011110111100010101010111010101;
12'b100010110101: dataB <= 32'b00001000000110101100010010011100;
12'b100010110110: dataB <= 32'b10010100110100110100001011010011;
12'b100010110111: dataB <= 32'b00000101011001100101101001111011;
12'b100010111000: dataB <= 32'b11100110001110011101010100110001;
12'b100010111001: dataB <= 32'b00001010011110101101011110111001;
12'b100010111010: dataB <= 32'b00001101011001111111101000010111;
12'b100010111011: dataB <= 32'b00000100111101011011011001011110;
12'b100010111100: dataB <= 32'b11011111010010000110100100110101;
12'b100010111101: dataB <= 32'b00001010101001111010101000001011;
12'b100010111110: dataB <= 32'b10010110000101101011000100001001;
12'b100010111111: dataB <= 32'b00000111100001100110001101110000;
12'b100011000000: dataB <= 32'b01011010101001110111101001011001;
12'b100011000001: dataB <= 32'b00001010000001101110010110001011;
12'b100011000010: dataB <= 32'b00000011001101010010000011100100;
12'b100011000011: dataB <= 32'b00000111010100101001011000011110;
12'b100011000100: dataB <= 32'b01111100110000111010101101010011;
12'b100011000101: dataB <= 32'b00000111101010101010101111100011;
12'b100011000110: dataB <= 32'b01011111000001011101010100010001;
12'b100011000111: dataB <= 32'b00000000110011101011110101001100;
12'b100011001000: dataB <= 32'b00101111100001010001010111100110;
12'b100011001001: dataB <= 32'b00000010001010010000110010111111;
12'b100011001010: dataB <= 32'b10101111010010001111001100011100;
12'b100011001011: dataB <= 32'b00000000110100010001001110010100;
12'b100011001100: dataB <= 32'b11111000100000101110100001110100;
12'b100011001101: dataB <= 32'b00001000000111101100010000111000;
12'b100011001110: dataB <= 32'b01010110111110010101110010101101;
12'b100011001111: dataB <= 32'b00001101000110101100010000101011;
12'b100011010000: dataB <= 32'b10100110011101111111100010010000;
12'b100011010001: dataB <= 32'b00001110110111011000101101110001;
12'b100011010010: dataB <= 32'b11101101011001010010110111101100;
12'b100011010011: dataB <= 32'b00000011000101010100001000011011;
12'b100011010100: dataB <= 32'b11011100000111001010100111000101;
12'b100011010101: dataB <= 32'b00000011011011011011100110000001;
12'b100011010110: dataB <= 32'b00110000110001010111100101110101;
12'b100011010111: dataB <= 32'b00001101000101111010101010011011;
12'b100011011000: dataB <= 32'b10010010111010100111100110001111;
12'b100011011001: dataB <= 32'b00000010101000101000110101110100;
12'b100011011010: dataB <= 32'b00010000101001110111100110011000;
12'b100011011011: dataB <= 32'b00001100101001010110000110011100;
12'b100011011100: dataB <= 32'b11000010101010101110100001001110;
12'b100011011101: dataB <= 32'b00000100010000101011011010001100;
12'b100011011110: dataB <= 32'b01111001011101100010011111001101;
12'b100011011111: dataB <= 32'b00000100110100001011000101000011;
12'b100011100000: dataB <= 32'b00100000001101110110011001111001;
12'b100011100001: dataB <= 32'b00001101110000111100110001111010;
12'b100011100010: dataB <= 32'b00111100111000011100000100010000;
12'b100011100011: dataB <= 32'b00001001111000011001001011001011;
12'b100011100100: dataB <= 32'b10001100010101100001010100100010;
12'b100011100101: dataB <= 32'b00000000110001001011001110000010;
12'b100011100110: dataB <= 32'b10001011011001100011011000101110;
12'b100011100111: dataB <= 32'b00001011001100011110000100010101;
12'b100011101000: dataB <= 32'b00101101001100110001011111001111;
12'b100011101001: dataB <= 32'b00001010110100100101000011100110;
12'b100011101010: dataB <= 32'b10010110100101110010111101001111;
12'b100011101011: dataB <= 32'b00000110010111100011011100100001;
12'b100011101100: dataB <= 32'b11011110110101000101010111010011;
12'b100011101101: dataB <= 32'b00001010011110000010101000011010;
12'b100011101110: dataB <= 32'b10100011100010001011110010100111;
12'b100011101111: dataB <= 32'b00000011110001011001001000010101;
12'b100011110000: dataB <= 32'b10111010111010100010100111100111;
12'b100011110001: dataB <= 32'b00001000000001110110011101100001;
12'b100011110010: dataB <= 32'b01000010101000100101000100110101;
12'b100011110011: dataB <= 32'b00001011101000100110010110110101;
12'b100011110100: dataB <= 32'b00010010101111101101100010101000;
12'b100011110101: dataB <= 32'b00001001000001011000000110111101;
12'b100011110110: dataB <= 32'b00101110111110001011000100100010;
12'b100011110111: dataB <= 32'b00000101001010111101001101000010;
12'b100011111000: dataB <= 32'b00010001001101110111101010011110;
12'b100011111001: dataB <= 32'b00001011010011111011011000111111;
12'b100011111010: dataB <= 32'b10110000101101011001101000101000;
12'b100011111011: dataB <= 32'b00001011001110100010101101010001;
12'b100011111100: dataB <= 32'b00001101000001010110001011111100;
12'b100011111101: dataB <= 32'b00000010001010110101010000011101;
12'b100011111110: dataB <= 32'b11000110101100101101010001010001;
12'b100011111111: dataB <= 32'b00000001110111000011000001001011;
12'b100100000000: dataB <= 32'b11100110110100001100001101111001;
12'b100100000001: dataB <= 32'b00000000110001000100111001110010;
12'b100100000010: dataB <= 32'b11100001001110011010111011100011;
12'b100100000011: dataB <= 32'b00001110001011010110001000111011;
12'b100100000100: dataB <= 32'b11101001100100011101011000011011;
12'b100100000101: dataB <= 32'b00001011101101111000111000001011;
12'b100100000110: dataB <= 32'b10011111010010110010101001001000;
12'b100100000111: dataB <= 32'b00001100010111010100111110100111;
12'b100100001000: dataB <= 32'b10001000111010110100001000101101;
12'b100100001001: dataB <= 32'b00000111110010010110111111010110;
12'b100100001010: dataB <= 32'b10011110111100001100110110110101;
12'b100100001011: dataB <= 32'b00001001000111110000010110011100;
12'b100100001100: dataB <= 32'b10010110110000110011101010110101;
12'b100100001101: dataB <= 32'b00000100111000100001101001111011;
12'b100100001110: dataB <= 32'b01101100010010010101010100101111;
12'b100100001111: dataB <= 32'b00001001011110101001100011001010;
12'b100100010000: dataB <= 32'b11001011010001100111100111110111;
12'b100100010001: dataB <= 32'b00000011111100011001011001001101;
12'b100100010010: dataB <= 32'b00011111010001110110100100010100;
12'b100100010011: dataB <= 32'b00001011001011111010110100001011;
12'b100100010100: dataB <= 32'b10011100000101110010110100101000;
12'b100100010101: dataB <= 32'b00001001000001101010010010000000;
12'b100100010110: dataB <= 32'b01011100100101011111101000011001;
12'b100100010111: dataB <= 32'b00001011100010110010011110001011;
12'b100100011000: dataB <= 32'b01000011000001100001110100100011;
12'b100100011001: dataB <= 32'b00000110110100100101011100010101;
12'b100100011010: dataB <= 32'b00111100111101000010001100110101;
12'b100100011011: dataB <= 32'b00001000001010101100110011100100;
12'b100100011100: dataB <= 32'b11011111000001010101000100010000;
12'b100100011101: dataB <= 32'b00000000110000100101110101001011;
12'b100100011110: dataB <= 32'b10101011101001100001001000100110;
12'b100100011111: dataB <= 32'b00000010101000010010101010101111;
12'b100100100000: dataB <= 32'b10101101010101111111001010111101;
12'b100100100001: dataB <= 32'b00000000110010001111001010001100;
12'b100100100010: dataB <= 32'b10111100101100011110000001010010;
12'b100100100011: dataB <= 32'b00001000100111110000010101010000;
12'b100100100100: dataB <= 32'b11010110111110001101110011001011;
12'b100100100101: dataB <= 32'b00001110001001110000010100110010;
12'b100100100110: dataB <= 32'b10101000100001101111100010001110;
12'b100100100111: dataB <= 32'b00001101111001011010101101111001;
12'b100100101000: dataB <= 32'b00101011011101011010101000001100;
12'b100100101001: dataB <= 32'b00000100100011011010000100100011;
12'b100100101010: dataB <= 32'b11100010000111010011001000100101;
12'b100100101011: dataB <= 32'b00000010011001010111100010001001;
12'b100100101100: dataB <= 32'b00110010111001000111000101010100;
12'b100100101101: dataB <= 32'b00001110001000111100110110011011;
12'b100100101110: dataB <= 32'b10010100110110001111100110101110;
12'b100100101111: dataB <= 32'b00000011100110101000111001110100;
12'b100100110000: dataB <= 32'b01010010100101011111100101110111;
12'b100100110001: dataB <= 32'b00001101001011011100000110010100;
12'b100100110010: dataB <= 32'b11000110100010011110100001001011;
12'b100100110011: dataB <= 32'b00000100001111101001011110001100;
12'b100100110100: dataB <= 32'b00110101101001101010011111010000;
12'b100100110101: dataB <= 32'b00000100010010001010111001000011;
12'b100100110110: dataB <= 32'b00100110010001100110001000111010;
12'b100100110111: dataB <= 32'b00001101010010111100111110000010;
12'b100100111000: dataB <= 32'b10111101000100011011010100001111;
12'b100100111001: dataB <= 32'b00001000111001010111000111010011;
12'b100100111010: dataB <= 32'b10010010001101110001000101100001;
12'b100100111011: dataB <= 32'b00000000101110001001000110001010;
12'b100100111100: dataB <= 32'b11001001010001101011001001001111;
12'b100100111101: dataB <= 32'b00001011001101100100000100001100;
12'b100100111110: dataB <= 32'b10101011010001001000111111010010;
12'b100100111111: dataB <= 32'b00001010010101100101000011010110;
12'b100101000000: dataB <= 32'b00011010100001111010111101010001;
12'b100101000001: dataB <= 32'b00000101010110100001011100110001;
12'b100101000010: dataB <= 32'b01011110110100111100110111010011;
12'b100101000011: dataB <= 32'b00001000111110000110100000100010;
12'b100101000100: dataB <= 32'b11011111100010001011110011100101;
12'b100101000101: dataB <= 32'b00000011101111010111000100001100;
12'b100101000110: dataB <= 32'b01111011000010101010111000101000;
12'b100101000111: dataB <= 32'b00001001000001111000100101110001;
12'b100101001000: dataB <= 32'b10000110100000100100010100010100;
12'b100101001001: dataB <= 32'b00001100001010101010011010100101;
12'b100101001010: dataB <= 32'b01010100101011100110000011100110;
12'b100101001011: dataB <= 32'b00001010100001011110000110110101;
12'b100101001100: dataB <= 32'b11101111000010010011000101100001;
12'b100101001101: dataB <= 32'b00000101101010111011011001010001;
12'b100101001110: dataB <= 32'b10001111001001011111101000111110;
12'b100101001111: dataB <= 32'b00001010110100111001100000101110;
12'b100101010000: dataB <= 32'b01110000110001101001101001001001;
12'b100101010001: dataB <= 32'b00001011010000100100101101100001;
12'b100101010010: dataB <= 32'b10001100111001000101111010111110;
12'b100101010011: dataB <= 32'b00000010101000110011011000010100;
12'b100101010100: dataB <= 32'b10001000100100101100110001001111;
12'b100101010101: dataB <= 32'b00000000110101000010110101001011;
12'b100101010110: dataB <= 32'b11101000111000001011011100111011;
12'b100101010111: dataB <= 32'b00000000101110000100101101111010;
12'b100101011000: dataB <= 32'b10011111001110100010111101000101;
12'b100101011001: dataB <= 32'b00001110101101011100000100111011;
12'b100101011010: dataB <= 32'b01100101100100010100110111011011;
12'b100101011011: dataB <= 32'b00001011101110111001000000001011;
12'b100101011100: dataB <= 32'b10011111010010111010111001101000;
12'b100101011101: dataB <= 32'b00001011011001010100111010001111;
12'b100101011110: dataB <= 32'b00001000110010110100011000101101;
12'b100101011111: dataB <= 32'b00000111110010010110111111000111;
12'b100101100000: dataB <= 32'b11011110111100001100000110010100;
12'b100101100001: dataB <= 32'b00001010000111110100011110010100;
12'b100101100010: dataB <= 32'b10010110101100111011001010010101;
12'b100101100011: dataB <= 32'b00000011110111011101101001111011;
12'b100101100100: dataB <= 32'b11110000010110001101100100101110;
12'b100101100101: dataB <= 32'b00000111111110100111100011010010;
12'b100101100110: dataB <= 32'b10001001001001001111010110110111;
12'b100101100111: dataB <= 32'b00000010111010010111010101000101;
12'b100101101000: dataB <= 32'b01011101010001100110010011110010;
12'b100101101001: dataB <= 32'b00001011101100111100111100010010;
12'b100101101010: dataB <= 32'b10100010000101111010110101100111;
12'b100101101011: dataB <= 32'b00001010100001110000010110011000;
12'b100101101100: dataB <= 32'b10011110100101000111010111111001;
12'b100101101101: dataB <= 32'b00001100100100110110100110010011;
12'b100101101110: dataB <= 32'b10000010110101110001110110000010;
12'b100101101111: dataB <= 32'b00000110010011100011011100001100;
12'b100101110000: dataB <= 32'b10111101001001010001111100010111;
12'b100101110001: dataB <= 32'b00001000101010101110110111100100;
12'b100101110010: dataB <= 32'b10011111000001001100110100001110;
12'b100101110011: dataB <= 32'b00000000101101100001111001001011;
12'b100101110100: dataB <= 32'b10100111101101111000111001100111;
12'b100101110101: dataB <= 32'b00000011000110010100100110010111;
12'b100101110110: dataB <= 32'b10101011011001100110111001011110;
12'b100101110111: dataB <= 32'b00000000101111001111000010001100;
12'b100101111000: dataB <= 32'b01111100110100010101100001001111;
12'b100101111001: dataB <= 32'b00001001100111110100011101101000;
12'b100101111010: dataB <= 32'b10010110111001111101110011101010;
12'b100101111011: dataB <= 32'b00001110101011110100011100111010;
12'b100101111100: dataB <= 32'b10101100100101010111010010101100;
12'b100101111101: dataB <= 32'b00001100111011011100101010001001;
12'b100101111110: dataB <= 32'b10101001100001100010011000101100;
12'b100101111111: dataB <= 32'b00000101100010100000000100101010;
12'b100110000000: dataB <= 32'b11101000000111010011101001100101;
12'b100110000001: dataB <= 32'b00000001010111010011011110011001;
12'b100110000010: dataB <= 32'b01110011000000101110100100110011;
12'b100110000011: dataB <= 32'b00001111001010111101000010100011;
12'b100110000100: dataB <= 32'b01010100110001110111100110101110;
12'b100110000101: dataB <= 32'b00000100100100101000111101101100;
12'b100110000110: dataB <= 32'b01010110100001000111010100110110;
12'b100110000111: dataB <= 32'b00001101001101100010000110010100;
12'b100110001000: dataB <= 32'b11001010010110001110110001101001;
12'b100110001001: dataB <= 32'b00000100101101100101100010000100;
12'b100110001010: dataB <= 32'b11110001110001111010001111010011;
12'b100110001011: dataB <= 32'b00000100010001001010110001001010;
12'b100110001100: dataB <= 32'b01101010010101010110000111111010;
12'b100110001101: dataB <= 32'b00001101010100111101001010010010;
12'b100110001110: dataB <= 32'b00111101010000100010110100101101;
12'b100110001111: dataB <= 32'b00000111111001010111000011010100;
12'b100110010000: dataB <= 32'b11010110001010001001000111000001;
12'b100110010001: dataB <= 32'b00000000101011001000111010010010;
12'b100110010010: dataB <= 32'b00000111001001110011001001001111;
12'b100110010011: dataB <= 32'b00001011101111101010000100001100;
12'b100110010100: dataB <= 32'b00101001010101011000101111010101;
12'b100110010101: dataB <= 32'b00001001110110100101000010111111;
12'b100110010110: dataB <= 32'b10011100100010000010111100110011;
12'b100110010111: dataB <= 32'b00000100110101011101011101000000;
12'b100110011000: dataB <= 32'b11100000110100111100010110110011;
12'b100110011001: dataB <= 32'b00000111011110001010010100110001;
12'b100110011010: dataB <= 32'b00011011100010001100000101000100;
12'b100110011011: dataB <= 32'b00000011101101010111000000001100;
12'b100110011100: dataB <= 32'b01111011001110110011001001001000;
12'b100110011101: dataB <= 32'b00001010100010111010110010000001;
12'b100110011110: dataB <= 32'b11001010010100011011110011110010;
12'b100110011111: dataB <= 32'b00001100101011101110011110011101;
12'b100110100000: dataB <= 32'b10010110100111010110100100100100;
12'b100110100001: dataB <= 32'b00001011100011100100000110101101;
12'b100110100010: dataB <= 32'b10101101001010011011010111000001;
12'b100110100011: dataB <= 32'b00000110101001111001100001011001;
12'b100110100100: dataB <= 32'b11001111000001000111010111011110;
12'b100110100101: dataB <= 32'b00001010010101110101101000011101;
12'b100110100110: dataB <= 32'b01110010111001111001101010001010;
12'b100110100111: dataB <= 32'b00001011010001100110110001110001;
12'b100110101000: dataB <= 32'b11001110110000111101011001011110;
12'b100110101001: dataB <= 32'b00000011000110101111011100010011;
12'b100110101010: dataB <= 32'b01001100011100100100010001001100;
12'b100110101011: dataB <= 32'b00000000110010000100101001001011;
12'b100110101100: dataB <= 32'b11101000111100001010111011111101;
12'b100110101101: dataB <= 32'b00000000101011000110100110000010;
12'b100110101110: dataB <= 32'b00011101001110101011001110000111;
12'b100110101111: dataB <= 32'b00001110110000100010000100111011;
12'b100110110000: dataB <= 32'b10100001100100010100000110011010;
12'b100110110001: dataB <= 32'b00001011110000110111001100010010;
12'b100110110010: dataB <= 32'b10011101010011000011011010001001;
12'b100110110011: dataB <= 32'b00001010011010010110110101110111;
12'b100110110100: dataB <= 32'b01001010101010110100101001001110;
12'b100110110101: dataB <= 32'b00000111110010010110111010110111;
12'b100110110110: dataB <= 32'b11011110111100001011010101110011;
12'b100110110111: dataB <= 32'b00001010101000110110101010001100;
12'b100110111000: dataB <= 32'b10011000101000111010101001010110;
12'b100110111001: dataB <= 32'b00000011010101011001100110000011;
12'b100110111010: dataB <= 32'b01110100011110000101100100101101;
12'b100110111011: dataB <= 32'b00000110011110100011100111010011;
12'b100110111100: dataB <= 32'b00001001000000111111000110010110;
12'b100110111101: dataB <= 32'b00000001110111010101010000111101;
12'b100110111110: dataB <= 32'b11011011001101010110000011110001;
12'b100110111111: dataB <= 32'b00001011101101111011001000011001;
12'b100111000000: dataB <= 32'b11101000000101111010110110100110;
12'b100111000001: dataB <= 32'b00001011100011110100011110101000;
12'b100111000010: dataB <= 32'b10100010100100110110110110111001;
12'b100111000011: dataB <= 32'b00001101100110111000101110010011;
12'b100111000100: dataB <= 32'b00000100101001111001110111100001;
12'b100111000101: dataB <= 32'b00000110010011011111100000001100;
12'b100111000110: dataB <= 32'b01111101010101100001101011011000;
12'b100111000111: dataB <= 32'b00001001001010101110111111011101;
12'b100111001000: dataB <= 32'b01011111000001001100100100001101;
12'b100111001001: dataB <= 32'b00000001001010011011110101010011;
12'b100111001010: dataB <= 32'b10100011101110001000111010000111;
12'b100111001011: dataB <= 32'b00000100000101011000100001111111;
12'b100111001100: dataB <= 32'b11101001011101010110101000011110;
12'b100111001101: dataB <= 32'b00000000101100001110111010000100;
12'b100111001110: dataB <= 32'b01111101000000001100110001001100;
12'b100111001111: dataB <= 32'b00001010101000110110100101111000;
12'b100111010000: dataB <= 32'b00011000110101110101110100001000;
12'b100111010001: dataB <= 32'b00001110101110110110100101000010;
12'b100111010010: dataB <= 32'b11101110101000111111000010101010;
12'b100111010011: dataB <= 32'b00001011111101011110101010011001;
12'b100111010100: dataB <= 32'b00100101100001101010011000101100;
12'b100111010101: dataB <= 32'b00000111000010100110000100110010;
12'b100111010110: dataB <= 32'b00101110001011010100011010100110;
12'b100111010111: dataB <= 32'b00000000110100010001011010101010;
12'b100111011000: dataB <= 32'b10110011000100011110000100110010;
12'b100111011001: dataB <= 32'b00001111001101111101001110100011;
12'b100111011010: dataB <= 32'b01010110101101011111100110101101;
12'b100111011011: dataB <= 32'b00000101100011101001000001101100;
12'b100111011100: dataB <= 32'b10011000011100110110110100010101;
12'b100111011101: dataB <= 32'b00001101101111101000000110010100;
12'b100111011110: dataB <= 32'b11001110001101111110110010100110;
12'b100111011111: dataB <= 32'b00000100101100100011100001111100;
12'b100111100000: dataB <= 32'b01101101110110000010001110110110;
12'b100111100001: dataB <= 32'b00000011101111001100101001010010;
12'b100111100010: dataB <= 32'b01101110011001001101100110111010;
12'b100111100011: dataB <= 32'b00001100110110111101010010011010;
12'b100111100100: dataB <= 32'b10111011011100101010010100101100;
12'b100111100101: dataB <= 32'b00000111011001010111000011010100;
12'b100111100110: dataB <= 32'b11011100001010011001011000100001;
12'b100111100111: dataB <= 32'b00000001001001001010110010011010;
12'b100111101000: dataB <= 32'b01000110111101110011001001001111;
12'b100111101001: dataB <= 32'b00001011110000101110001100001011;
12'b100111101010: dataB <= 32'b10100111011001110000101110010111;
12'b100111101011: dataB <= 32'b00001001010110100011000110101111;
12'b100111101100: dataB <= 32'b01100000011110001010111100010101;
12'b100111101101: dataB <= 32'b00000100010011011011011101011000;
12'b100111101110: dataB <= 32'b01100000110100111100000110010010;
12'b100111101111: dataB <= 32'b00000101111110001110001101000001;
12'b100111110000: dataB <= 32'b01011001011110001100000110000011;
12'b100111110001: dataB <= 32'b00000100001100010111000000001011;
12'b100111110010: dataB <= 32'b01111001010110110011011010001001;
12'b100111110011: dataB <= 32'b00001100000011111100111110010001;
12'b100111110100: dataB <= 32'b11001110001100100011010011110001;
12'b100111110101: dataB <= 32'b00001101001101110000100110010101;
12'b100111110110: dataB <= 32'b11011010100010111111000101100011;
12'b100111110111: dataB <= 32'b00001101000101101010001010100101;
12'b100111111000: dataB <= 32'b01101101001110011011101000100001;
12'b100111111001: dataB <= 32'b00000111001000110101101001101001;
12'b100111111010: dataB <= 32'b01001110111000110110110101111110;
12'b100111111011: dataB <= 32'b00001001110110101111110000001101;
12'b100111111100: dataB <= 32'b01110011000010001001101010101010;
12'b100111111101: dataB <= 32'b00001010110010100110110010001001;
12'b100111111110: dataB <= 32'b00001110101100110100110111111110;
12'b100111111111: dataB <= 32'b00000100000101101101100100010011;
12'b101000000000: dataB <= 32'b00010000010100100011110001101010;
12'b101000000001: dataB <= 32'b00000000101111000110011101010011;
12'b101000000010: dataB <= 32'b11101000111100011010001010011110;
12'b101000000011: dataB <= 32'b00000001001000001010011010001010;
12'b101000000100: dataB <= 32'b10011101001110101011101110101001;
12'b101000000101: dataB <= 32'b00001110110011101000001001000010;
12'b101000000110: dataB <= 32'b11011101100100010011100101011010;
12'b101000000111: dataB <= 32'b00001011110001110101010100011001;
12'b101000001000: dataB <= 32'b10011011001111000011101011001010;
12'b101000001001: dataB <= 32'b00001001011011010110110001011111;
12'b101000001010: dataB <= 32'b10001110100010101100111001001110;
12'b101000001011: dataB <= 32'b00000111010001011000110110011111;
12'b101000001100: dataB <= 32'b11011110111100010010100101010010;
12'b101000001101: dataB <= 32'b00001011001001111000110010001100;
12'b101000001110: dataB <= 32'b10011100101001001010011000110111;
12'b101000001111: dataB <= 32'b00000010110011010101100010000011;
12'b101000010000: dataB <= 32'b11110110100101110101100101001100;
12'b101000010001: dataB <= 32'b00000100111101011111100111011011;
12'b101000010010: dataB <= 32'b10001000111000101110100101110101;
12'b101000010011: dataB <= 32'b00000000110101010011001100110100;
12'b101000010100: dataB <= 32'b00011001001101000101110011101111;
12'b101000010101: dataB <= 32'b00001100001111111011010100101001;
12'b101000010110: dataB <= 32'b01101110001010000010110111100101;
12'b101000010111: dataB <= 32'b00001101000100110110100111000001;
12'b101000011000: dataB <= 32'b11100100101000100110010101111000;
12'b101000011001: dataB <= 32'b00001110101000111010111010010011;
12'b101000011010: dataB <= 32'b01000110011110001001111000100001;
12'b101000011011: dataB <= 32'b00000101110010011101011100001011;
12'b101000011100: dataB <= 32'b11111001011101110001101010111001;
12'b101000011101: dataB <= 32'b00001001101011101111000011010101;
12'b101000011110: dataB <= 32'b00011111000001001100010100101011;
12'b101000011111: dataB <= 32'b00000001100111010101110101010011;
12'b101000100000: dataB <= 32'b10011111101110011001001011001000;
12'b101000100001: dataB <= 32'b00000101100011011010100001100111;
12'b101000100010: dataB <= 32'b11100101100001000110010110111110;
12'b101000100011: dataB <= 32'b00000001001001001110110101111100;
12'b101000100100: dataB <= 32'b01111101001100001100000001101010;
12'b101000100101: dataB <= 32'b00001011001001111000110010010000;
12'b101000100110: dataB <= 32'b11011000110001100101110101000111;
12'b101000100111: dataB <= 32'b00001110110001111000110001010001;
12'b101000101000: dataB <= 32'b00110000110000101110100011101000;
12'b101000101001: dataB <= 32'b00001010011110100000101010100010;
12'b101000101010: dataB <= 32'b10100001100101110010011001001101;
12'b101000101011: dataB <= 32'b00001000100010101010001001000001;
12'b101000101100: dataB <= 32'b01110010010011010100111011000111;
12'b101000101101: dataB <= 32'b00000000110001001111010010110010;
12'b101000101110: dataB <= 32'b11110001001100010101100100110001;
12'b101000101111: dataB <= 32'b00001111010000111011010110101011;
12'b101000110000: dataB <= 32'b00011000101001000111010111001101;
12'b101000110001: dataB <= 32'b00000111000010101001000101101100;
12'b101000110010: dataB <= 32'b10011100011100100110010011110011;
12'b101000110011: dataB <= 32'b00001101110001101110001010001100;
12'b101000110100: dataB <= 32'b11010010001001101110110011100101;
12'b101000110101: dataB <= 32'b00000101001011011111100001110100;
12'b101000110110: dataB <= 32'b00100111111010010010011101111001;
12'b101000110111: dataB <= 32'b00000100001110001110100101011010;
12'b101000111000: dataB <= 32'b10110010100001000101010101111001;
12'b101000111001: dataB <= 32'b00001011111000111001011110100010;
12'b101000111010: dataB <= 32'b00110111100100111001110101001011;
12'b101000111011: dataB <= 32'b00000110011000010110111111001101;
12'b101000111100: dataB <= 32'b00100010001010101001101010000001;
12'b101000111101: dataB <= 32'b00000010000110001100101010100011;
12'b101000111110: dataB <= 32'b11000110110101111010111001010000;
12'b101000111111: dataB <= 32'b00001011010010110100010000001010;
12'b101001000000: dataB <= 32'b10100101011010001000101101111010;
12'b101001000001: dataB <= 32'b00001000110110100011000110010111;
12'b101001000010: dataB <= 32'b01100010100010001011001011110111;
12'b101001000011: dataB <= 32'b00000100010010010111011001110000;
12'b101001000100: dataB <= 32'b00100010110100111011100110010010;
12'b101001000101: dataB <= 32'b00000100011101010010001001010001;
12'b101001000110: dataB <= 32'b11010101011010001100000111100010;
12'b101001000111: dataB <= 32'b00000100101010010110111100001010;
12'b101001001000: dataB <= 32'b10110101100010110011101010101010;
12'b101001001001: dataB <= 32'b00001101000101111101000110100001;
12'b101001001010: dataB <= 32'b00010010001000101010100011101111;
12'b101001001011: dataB <= 32'b00001101001111110010101010000110;
12'b101001001100: dataB <= 32'b00011100100010101111100111000010;
12'b101001001101: dataB <= 32'b00001110000111110000001110010110;
12'b101001001110: dataB <= 32'b01101011010010011011101010000001;
12'b101001001111: dataB <= 32'b00000111101000101111110001111001;
12'b101001010000: dataB <= 32'b10001110110100100110010100011101;
12'b101001010001: dataB <= 32'b00001001010110101011111000001100;
12'b101001010010: dataB <= 32'b01110011001010011001101011001100;
12'b101001010011: dataB <= 32'b00001010110011101000110110011001;
12'b101001010100: dataB <= 32'b10010000100100110100010110011110;
12'b101001010101: dataB <= 32'b00000101100011101001101000011010;
12'b101001010110: dataB <= 32'b11010100010000100011010010100111;
12'b101001010111: dataB <= 32'b00000000101100001010010101011010;
12'b101001011000: dataB <= 32'b00101001000000100001101000111110;
12'b101001011001: dataB <= 32'b00000010000110001110010110001011;
12'b101001011010: dataB <= 32'b01011011001010110011111111001100;
12'b101001011011: dataB <= 32'b00001110010101101100001101001010;
12'b101001011100: dataB <= 32'b01011001100100011010110100011000;
12'b101001011101: dataB <= 32'b00001011110011110011011100101001;
12'b101001011110: dataB <= 32'b01011001001111000100001011101011;
12'b101001011111: dataB <= 32'b00001000011011011000101101000111;
12'b101001100000: dataB <= 32'b10010000011010100101001001001111;
12'b101001100001: dataB <= 32'b00000111010001011000110010000111;
12'b101001100010: dataB <= 32'b00011110111100011001110101010001;
12'b101001100011: dataB <= 32'b00001100001011111010111110000101;
12'b101001100100: dataB <= 32'b10011110100101010010001000010111;
12'b101001100101: dataB <= 32'b00000010010001010001011110000011;
12'b101001100110: dataB <= 32'b01111000110001101101010101101011;
12'b101001100111: dataB <= 32'b00000011011011011011100111011100;
12'b101001101000: dataB <= 32'b00001010101100011101110101010100;
12'b101001101001: dataB <= 32'b00000000110010010011001000101100;
12'b101001101010: dataB <= 32'b11011001001000111101010011101101;
12'b101001101011: dataB <= 32'b00001100010001110111011101000000;
12'b101001101100: dataB <= 32'b10110010010010001010111000100101;
12'b101001101101: dataB <= 32'b00001110000111111000101111010001;
12'b101001101110: dataB <= 32'b11100110101000010101100100110111;
12'b101001101111: dataB <= 32'b00001111001011111011000010010011;
12'b101001110000: dataB <= 32'b10001010010110011001111010000010;
12'b101001110001: dataB <= 32'b00000101110001011001011100010010;
12'b101001110010: dataB <= 32'b01110101101010000001011001111010;
12'b101001110011: dataB <= 32'b00001010001100101111001011000110;
12'b101001110100: dataB <= 32'b11011111000001000011110101001010;
12'b101001110101: dataB <= 32'b00000010100101010001101101011010;
12'b101001110110: dataB <= 32'b01011011101110101001011011101010;
12'b101001110111: dataB <= 32'b00000110100011011110100001001111;
12'b101001111000: dataB <= 32'b11100001100000110101110101011101;
12'b101001111001: dataB <= 32'b00000010000111010000101101111100;
12'b101001111010: dataB <= 32'b10111011011000001011010010101000;
12'b101001111011: dataB <= 32'b00001011101011111000111010101000;
12'b101001111100: dataB <= 32'b10011010110001011101100110000110;
12'b101001111101: dataB <= 32'b00001110110011111000111001100001;
12'b101001111110: dataB <= 32'b01110000111000011110000100100110;
12'b101001111111: dataB <= 32'b00001000111110100010101010110010;
12'b101010000000: dataB <= 32'b01011101100110000010001001001101;
12'b101010000001: dataB <= 32'b00001001100010110000001101001001;
12'b101010000010: dataB <= 32'b11110110011011001101011100001001;
12'b101010000011: dataB <= 32'b00000000101110001101001010111010;
12'b101010000100: dataB <= 32'b00101111010100001100110100001111;
12'b101010000101: dataB <= 32'b00001111010011111001100010101100;
12'b101010000110: dataB <= 32'b00011010101000110110110111001101;
12'b101010000111: dataB <= 32'b00001000000010101001001001101100;
12'b101010001000: dataB <= 32'b10100000011000010101100011110001;
12'b101010001001: dataB <= 32'b00001101010011110010010010001100;
12'b101010001010: dataB <= 32'b11011000000101011110100100100011;
12'b101010001011: dataB <= 32'b00000101101010011011100001110100;
12'b101010001100: dataB <= 32'b00100001111010011010011101011011;
12'b101010001101: dataB <= 32'b00000100001100010010011101101010;
12'b101010001110: dataB <= 32'b11110100100100111100110100111000;
12'b101010001111: dataB <= 32'b00001010111001110111100110101010;
12'b101010010000: dataB <= 32'b10110011101101000001010101101010;
12'b101010010001: dataB <= 32'b00000101010111010110111011000101;
12'b101010010010: dataB <= 32'b01100110001010111001111011100010;
12'b101010010011: dataB <= 32'b00000011000100001110100010100011;
12'b101010010100: dataB <= 32'b00001000101110000010111001010000;
12'b101010010101: dataB <= 32'b00001011010011111000011100011010;
12'b101010010110: dataB <= 32'b10100001011010011000101100011100;
12'b101010010111: dataB <= 32'b00000111110111100011000101111111;
12'b101010011000: dataB <= 32'b01100110100010010011001010111000;
12'b101010011001: dataB <= 32'b00000100010000010101010110001000;
12'b101010011010: dataB <= 32'b11100010110100111011000110010001;
12'b101010011011: dataB <= 32'b00000011011011011000000101100000;
12'b101010011100: dataB <= 32'b00010011010110001100001000100010;
12'b101010011101: dataB <= 32'b00000101001001010110111000011010;
12'b101010011110: dataB <= 32'b11110011101010111100001011001011;
12'b101010011111: dataB <= 32'b00001110000111111011010010110001;
12'b101010100000: dataB <= 32'b00011000000100110010000011101101;
12'b101010100001: dataB <= 32'b00001101010010110100110001110110;
12'b101010100010: dataB <= 32'b00100000011110010111101000000010;
12'b101010100011: dataB <= 32'b00001110101001110100010110000110;
12'b101010100100: dataB <= 32'b01101001010110011011111011100010;
12'b101010100101: dataB <= 32'b00001000101000101011111010010001;
12'b101010100110: dataB <= 32'b11010000101100010101100011011011;
12'b101010100111: dataB <= 32'b00001000010110100101111000001011;
12'b101010101000: dataB <= 32'b10110001010010101001111011001101;
12'b101010101001: dataB <= 32'b00001010010100101000111010101001;
12'b101010101010: dataB <= 32'b00010100100000101011110100111101;
12'b101010101011: dataB <= 32'b00000110100011100101101000101010;
12'b101010101100: dataB <= 32'b10011000001100101010110011000101;
12'b101010101101: dataB <= 32'b00000001001001001110001101100010;
12'b101010101110: dataB <= 32'b00101001000100110001000111011110;
12'b101010101111: dataB <= 32'b00000011000100010010001110010011;
12'b101010110000: dataB <= 32'b00011011001010110100001111001111;
12'b101010110001: dataB <= 32'b00001101010111110000010101011010;
12'b101010110010: dataB <= 32'b11010101100000100010010011010110;
12'b101010110011: dataB <= 32'b00001011010100101111100100111000;
12'b101010110100: dataB <= 32'b11011001001011000100101011101101;
12'b101010110101: dataB <= 32'b00000111011011011010101100110110;
12'b101010110110: dataB <= 32'b10010100010110011101011001001111;
12'b101010110111: dataB <= 32'b00000111010001011010110001101111;
12'b101010111000: dataB <= 32'b00011110111100101001010101010000;
12'b101010111001: dataB <= 32'b00001100001101111011000101111101;
12'b101010111010: dataB <= 32'b10100000100101100001110111010111;
12'b101010111011: dataB <= 32'b00000010001111001111010110000011;
12'b101010111100: dataB <= 32'b11111000111001100101010110001010;
12'b101010111101: dataB <= 32'b00000010011010010111100011010100;
12'b101010111110: dataB <= 32'b10001100100100001101010100110011;
12'b101010111111: dataB <= 32'b00000000101111010011000000101011;
endcase
end
assign doA = dataA;
assign doB = dataB;
endmodule
