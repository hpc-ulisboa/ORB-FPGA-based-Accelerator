module rams_sp_rom0_4_sec (clk, enA, enB, addrA, addrB, doA, doB);
input clk;
input enA, enB;
input [10:0] addrA, addrB;
output [31:0] doA, doB;
(*rom_style = "block" *) reg [1375:0] dataA, dataB;
always @(posedge clk)
begin
if (enA)
case(addrA)
11'b00000000000: dataA <= 32'b00100101001110110101110111011000;
11'b00000000001: dataA <= 32'b00001000000111101100001100011110;
11'b00000000010: dataA <= 32'b10000110011101011011100010101111;
11'b00000000011: dataA <= 32'b00000010100100010100001100110001;
11'b00000000100: dataA <= 32'b01010100110111000111001100010101;
11'b00000000101: dataA <= 32'b00000101000010011110001001111011;
11'b00000000110: dataA <= 32'b10001101101100111011010001001100;
11'b00000000111: dataA <= 32'b00001000110100101111001001011111;
11'b00000001000: dataA <= 32'b10110010010000101100001101001011;
11'b00000001001: dataA <= 32'b00000110001011100010100011000001;
11'b00000001010: dataA <= 32'b00100001000010000101110101110110;
11'b00000001011: dataA <= 32'b00000011011011111001011001011101;
11'b00000001100: dataA <= 32'b01110111000100100010110100101001;
11'b00000001101: dataA <= 32'b00000001110011010001000111110101;
11'b00000001110: dataA <= 32'b00110000111011000110001111010100;
11'b00000001111: dataA <= 32'b00000100011100011001011110011100;
11'b00000010000: dataA <= 32'b11101010000101111111100100111011;
11'b00000010001: dataA <= 32'b00000101001000011010001100001010;
11'b00000010010: dataA <= 32'b00011001001010110100110011010100;
11'b00000010011: dataA <= 32'b00001001000010011010001100110101;
11'b00000010100: dataA <= 32'b10011010011111001110110011110111;
11'b00000010101: dataA <= 32'b00001111001101010100111101000010;
11'b00000010110: dataA <= 32'b11110011000001000100000110101101;
11'b00000010111: dataA <= 32'b00000001001101000100100000110101;
11'b00000011000: dataA <= 32'b00001010010110100001100100001000;
11'b00000011001: dataA <= 32'b00000111111110100111100101010010;
11'b00000011010: dataA <= 32'b10101000011110100111101000010111;
11'b00000011011: dataA <= 32'b00001000100001101110001010000010;
11'b00000011100: dataA <= 32'b10010101001111100110000110110001;
11'b00000011101: dataA <= 32'b00000001010000100100101110000100;
11'b00000011110: dataA <= 32'b10001101000011000111001001011000;
11'b00000011111: dataA <= 32'b00001001000101000110011110010011;
11'b00000100000: dataA <= 32'b01000011010011010100110010010111;
11'b00000100001: dataA <= 32'b00000101010101110001000110011100;
11'b00000100010: dataA <= 32'b11111100111001001011011101000100;
11'b00000100011: dataA <= 32'b00000110110111010001011101000100;
11'b00000100100: dataA <= 32'b10010000011010100110001100110101;
11'b00000100101: dataA <= 32'b00001100001001110000010001010010;
11'b00000100110: dataA <= 32'b10110100010100110110000101010101;
11'b00000100111: dataA <= 32'b00001100010100011101010010101001;
11'b00000101000: dataA <= 32'b11000100110100110010010001001010;
11'b00000101001: dataA <= 32'b00000010111010010011100101101010;
11'b00000101010: dataA <= 32'b01011001101101011011111000001101;
11'b00000101011: dataA <= 32'b00001001001001001010010001001111;
11'b00000101100: dataA <= 32'b11101100111000010011011101100101;
11'b00000101101: dataA <= 32'b00001011101111100010111011110011;
11'b00000101110: dataA <= 32'b11010000110101100011011011101001;
11'b00000101111: dataA <= 32'b00001000110111101101010000001011;
11'b00000110000: dataA <= 32'b00011010111001101110001000110011;
11'b00000110001: dataA <= 32'b00001110011000000011010000011101;
11'b00000110010: dataA <= 32'b01101101010110000011100001001111;
11'b00000110011: dataA <= 32'b00000101010110011101010001001111;
11'b00000110100: dataA <= 32'b10110010011001111010000101001001;
11'b00000110101: dataA <= 32'b00000011000100100110001000110010;
11'b00000110110: dataA <= 32'b00000011010001001110100111011000;
11'b00000110111: dataA <= 32'b00001000000101010110010111000100;
11'b00000111000: dataA <= 32'b10001111000011110011000001010000;
11'b00000111001: dataA <= 32'b00000100000010001000011011000011;
11'b00000111010: dataA <= 32'b11101010101001111011000001001010;
11'b00000111011: dataA <= 32'b00000100001111111010100100101011;
11'b00000111100: dataA <= 32'b10011001011111000111001110011000;
11'b00000111101: dataA <= 32'b00001011001110111100110010000111;
11'b00000111110: dataA <= 32'b11100110011100110010110110001001;
11'b00000111111: dataA <= 32'b00001010001011011100101100110010;
11'b00001000000: dataA <= 32'b11010011011010000110101111010101;
11'b00001000001: dataA <= 32'b00000001110011110100110001001110;
11'b00001000010: dataA <= 32'b00000111010001100110100011011001;
11'b00001000011: dataA <= 32'b00000101011110001001100101010101;
11'b00001000100: dataA <= 32'b01100010101100101110101111010000;
11'b00001000101: dataA <= 32'b00000010111010001001011101100011;
11'b00001000110: dataA <= 32'b01100101001001111010010111000001;
11'b00001000111: dataA <= 32'b00001011000100001000100001000101;
11'b00001001000: dataA <= 32'b01110011010001010111001011111000;
11'b00001001001: dataA <= 32'b00001001101001110000011100100110;
11'b00001001010: dataA <= 32'b00100101001110001001110110001000;
11'b00001001011: dataA <= 32'b00001101110000010111001011100110;
11'b00001001100: dataA <= 32'b00001011011010101010110111101101;
11'b00001001101: dataA <= 32'b00001000110001011001001011110100;
11'b00001001110: dataA <= 32'b00011111000000110110111000110101;
11'b00001001111: dataA <= 32'b00000110000111100000001010100100;
11'b00001010000: dataA <= 32'b11010011000000111101001011110000;
11'b00001010001: dataA <= 32'b00001000011011101101011101110011;
11'b00001010010: dataA <= 32'b01011010001110101100100101010100;
11'b00001010011: dataA <= 32'b00001101111010110001001110010001;
11'b00001010100: dataA <= 32'b10010101101010110111011010010110;
11'b00001010101: dataA <= 32'b00001000011110100011011001111110;
11'b00001010110: dataA <= 32'b00100111001011001101001000111000;
11'b00001010111: dataA <= 32'b00000110101000100010000101000111;
11'b00001011000: dataA <= 32'b11000010110101011100000011010011;
11'b00001011001: dataA <= 32'b00000001001001001100011000011010;
11'b00001011010: dataA <= 32'b01010010111111100110001100110001;
11'b00001011011: dataA <= 32'b00000010100101010100010001110011;
11'b00001011100: dataA <= 32'b10010111111000111100010000110010;
11'b00001011101: dataA <= 32'b00001001110011110000111110001111;
11'b00001011110: dataA <= 32'b11100110000100111101001100001000;
11'b00001011111: dataA <= 32'b00000101001101011100100010011000;
11'b00001100000: dataA <= 32'b10100001000010011101100110110111;
11'b00001100001: dataA <= 32'b00000101111110111101000101110101;
11'b00001100010: dataA <= 32'b11110110110100011011110011101100;
11'b00001100011: dataA <= 32'b00000010111000010011010011110011;
11'b00001100100: dataA <= 32'b11101110101011011101001111001110;
11'b00001100101: dataA <= 32'b00000110111110011111100010011011;
11'b00001100110: dataA <= 32'b01011110000110100111100111011101;
11'b00001100111: dataA <= 32'b00000100001011010000010100001100;
11'b00001101000: dataA <= 32'b00011011001110111100000100111000;
11'b00001101001: dataA <= 32'b00000110000010010000010101001110;
11'b00001101010: dataA <= 32'b01010100100111101101110101111010;
11'b00001101011: dataA <= 32'b00001110000111010101000100111011;
11'b00001101100: dataA <= 32'b10110000110001001100110110001110;
11'b00001101101: dataA <= 32'b00000001010011000010111001001110;
11'b00001101110: dataA <= 32'b11000100101001111001010011001011;
11'b00001101111: dataA <= 32'b00001010111101101111011101000010;
11'b00001110000: dataA <= 32'b11100010011011001110111001110110;
11'b00001110001: dataA <= 32'b00000110000001100010000101110010;
11'b00001110010: dataA <= 32'b10011001010011110100100111010010;
11'b00001110011: dataA <= 32'b00000010010101100000101110001100;
11'b00001110100: dataA <= 32'b01001111010011100110001010110110;
11'b00001110101: dataA <= 32'b00000111000100000010110110001011;
11'b00001110110: dataA <= 32'b11001001100111011011110011111011;
11'b00001110111: dataA <= 32'b00000110110110110000111010011011;
11'b00001111000: dataA <= 32'b10111000100001000100001010100001;
11'b00001111001: dataA <= 32'b00001000011000010111100101010101;
11'b00001111010: dataA <= 32'b01001010100110111101011101010001;
11'b00001111011: dataA <= 32'b00001010100110100110000101001011;
11'b00001111100: dataA <= 32'b01101010001001010110110110110110;
11'b00001111101: dataA <= 32'b00001100110001100001010010001001;
11'b00001111110: dataA <= 32'b00000101001100100011010000101111;
11'b00001111111: dataA <= 32'b00000101011101011011101101011011;
11'b00010000000: dataA <= 32'b10100011110001100100010111101101;
11'b00010000001: dataA <= 32'b00000111101000000100100101111111;
11'b00010000010: dataA <= 32'b01101010110000010100111011000010;
11'b00010000011: dataA <= 32'b00001011001100100010111011101010;
11'b00010000100: dataA <= 32'b01001111000001011011111010000110;
11'b00010000101: dataA <= 32'b00001010010110101111001000010101;
11'b00010000110: dataA <= 32'b00011010111110001110001001110010;
11'b00010000111: dataA <= 32'b00001111010010001001100100110110;
11'b00010001000: dataA <= 32'b10110001001110000011100001110100;
11'b00010001001: dataA <= 32'b00000110011000100001010001111111;
11'b00010001010: dataA <= 32'b10101000001101100010010100001100;
11'b00010001011: dataA <= 32'b00000001001000011010000100101011;
11'b00010001100: dataA <= 32'b01001001100101110110111000111000;
11'b00010001101: dataA <= 32'b00000110000110010000011110111011;
11'b00010001110: dataA <= 32'b10010001001111011001100010010101;
11'b00010001111: dataA <= 32'b00000010000110000010101110111010;
11'b00010010000: dataA <= 32'b11100100100101101011000000101111;
11'b00010010001: dataA <= 32'b00000100110010110010010000110100;
11'b00010010010: dataA <= 32'b01011111100011100110001111010010;
11'b00010010011: dataA <= 32'b00001010101100110110011010110111;
11'b00010010100: dataA <= 32'b00011110011000110011110101001011;
11'b00010010101: dataA <= 32'b00001000101001011000110000101100;
11'b00010010110: dataA <= 32'b01011001100010100110001111001111;
11'b00010010111: dataA <= 32'b00000010111000110000100101110111;
11'b00010011000: dataA <= 32'b01001101100010000110110101111100;
11'b00010011001: dataA <= 32'b00001000011110010011110101100101;
11'b00010011010: dataA <= 32'b11011110101101001111011110101010;
11'b00010011011: dataA <= 32'b00000101011101001111101101011011;
11'b00010011100: dataA <= 32'b11100111000101101010100100000011;
11'b00010011101: dataA <= 32'b00001000100010000100110101011101;
11'b00010011110: dataA <= 32'b01110011000001111111011101010100;
11'b00010011111: dataA <= 32'b00001000001000101000010001000111;
11'b00010100000: dataA <= 32'b10100111001001110001110100101010;
11'b00010100001: dataA <= 32'b00001101001100011001010011110100;
11'b00010100010: dataA <= 32'b11010011100110011010100111001101;
11'b00010100011: dataA <= 32'b00001000110001011011001111110010;
11'b00010100100: dataA <= 32'b10011111000001011111101001110100;
11'b00010100101: dataA <= 32'b00000100101001010110001110011011;
11'b00010100110: dataA <= 32'b11010101001001010101111011001101;
11'b00010100111: dataA <= 32'b00001010011010110011010001110011;
11'b00010101000: dataA <= 32'b00010000010110110100000110010101;
11'b00010101001: dataA <= 32'b00001111010101110010111101110001;
11'b00010101010: dataA <= 32'b01011111101111011110011011010100;
11'b00010101011: dataA <= 32'b00001011011101100111010110011110;
11'b00010101100: dataA <= 32'b10101001000011010100001010010110;
11'b00010101101: dataA <= 32'b00000101001001010110001001101111;
11'b00010101110: dataA <= 32'b00000011001001100100100100010111;
11'b00010101111: dataA <= 32'b00000000101111000110101100010100;
11'b00010110000: dataA <= 32'b10010011000111110100111100101110;
11'b00010110001: dataA <= 32'b00000001001010001100011101101011;
11'b00010110010: dataA <= 32'b01100011111001000101000001110111;
11'b00010110011: dataA <= 32'b00001010010001101110110010111111;
11'b00010110100: dataA <= 32'b11011100000101001101111010000101;
11'b00010110101: dataA <= 32'b00000101001111010110100101110000;
11'b00010110110: dataA <= 32'b10100001000010101101001000010111;
11'b00010110111: dataA <= 32'b00001000111110111010101110000101;
11'b00010111000: dataA <= 32'b01110010100100100101000011001111;
11'b00010111001: dataA <= 32'b00000100111011010111011011101010;
11'b00010111010: dataA <= 32'b10101010100011100011111110101000;
11'b00010111011: dataA <= 32'b00001001111110100111100010010011;
11'b00010111100: dataA <= 32'b11010010001011001110111001111101;
11'b00010111101: dataA <= 32'b00000011101110001010100000010101;
11'b00010111110: dataA <= 32'b01011111010010111011010110011001;
11'b00010111111: dataA <= 32'b00000011100100001010100001100110;
11'b00011000000: dataA <= 32'b01001110101111110100010111111011;
11'b00011000001: dataA <= 32'b00001100000011010111001100110100;
11'b00011000010: dataA <= 32'b11101100100101011101010110001111;
11'b00011000011: dataA <= 32'b00000010011000000011010001110110;
11'b00011000100: dataA <= 32'b10000010111101011001100010101111;
11'b00011000101: dataA <= 32'b00001101011010110011001100111011;
11'b00011000110: dataA <= 32'b00011010011111101101101010110100;
11'b00011000111: dataA <= 32'b00000011000100010110000101100011;
11'b00011001000: dataA <= 32'b01011101011011110011010111110011;
11'b00011001001: dataA <= 32'b00000011111001011100101110010100;
11'b00011001010: dataA <= 32'b00010101011011110100111100010100;
11'b00011001011: dataA <= 32'b00000101000110000011001010000011;
11'b00011001100: dataA <= 32'b10010011110111010010110110011101;
11'b00011001101: dataA <= 32'b00000111110111101100101110011011;
11'b00011001110: dataA <= 32'b11110010010001001100100111100001;
11'b00011001111: dataA <= 32'b00001001110111011111101001101101;
11'b00011010000: dataA <= 32'b11001000111011001100101101001101;
11'b00011010001: dataA <= 32'b00001000100100011010000101000011;
11'b00011010010: dataA <= 32'b01100000000101110111000111110111;
11'b00011010011: dataA <= 32'b00001100001101100101001101101001;
11'b00011010100: dataA <= 32'b10001001100000100100100001010101;
11'b00011010101: dataA <= 32'b00001000011110100101101101010011;
11'b00011010110: dataA <= 32'b10101011101101100100100111001110;
11'b00011010111: dataA <= 32'b00000110101001000010111110101111;
11'b00011011000: dataA <= 32'b00100110101000100110001000000001;
11'b00011011001: dataA <= 32'b00001010001010100000110111001001;
11'b00011011010: dataA <= 32'b10010001001101011100001000000101;
11'b00011011011: dataA <= 32'b00001011010100101110111100101110;
11'b00011011100: dataA <= 32'b11011011000010100101111001110001;
11'b00011011101: dataA <= 32'b00001111001101010011110101010110;
11'b00011011110: dataA <= 32'b10110000111101111011100011011001;
11'b00011011111: dataA <= 32'b00001000011000100101001110101111;
11'b00011100000: dataA <= 32'b10011110001001010010110011101111;
11'b00011100001: dataA <= 32'b00000000101110010000001100101100;
11'b00011100010: dataA <= 32'b10010011110110011110111010010110;
11'b00011100011: dataA <= 32'b00000100100111001010101110110010;
11'b00011100100: dataA <= 32'b00010101011010111000110011111001;
11'b00011100101: dataA <= 32'b00000000101100000011000110101010;
11'b00011100110: dataA <= 32'b10100000100001100011010001010101;
11'b00011100111: dataA <= 32'b00000101010100101000000100111101;
11'b00011101000: dataA <= 32'b01100111100011110100111111001101;
11'b00011101001: dataA <= 32'b00001001101010101110001111011110;
11'b00011101010: dataA <= 32'b00011000011100110100110100101101;
11'b00011101011: dataA <= 32'b00000111101001010110111000110101;
11'b00011101100: dataA <= 32'b01011111100110111101101110101001;
11'b00011101101: dataA <= 32'b00000100111011101010011010011111;
11'b00011101110: dataA <= 32'b10010101101110100110101000011101;
11'b00011101111: dataA <= 32'b00001011011101011101111001111101;
11'b00011110000: dataA <= 32'b00011010110001111111101101000101;
11'b00011110001: dataA <= 32'b00000111111110011001110101011100;
11'b00011110010: dataA <= 32'b00100111000001011010110010000110;
11'b00011110011: dataA <= 32'b00000110000010000101001001110110;
11'b00011110100: dataA <= 32'b10110010110010100111001101110000;
11'b00011110101: dataA <= 32'b00000110101000011110001101110111;
11'b00011110110: dataA <= 32'b01101001000001011010010100001101;
11'b00011110111: dataA <= 32'b00001100001000011101010111110011;
11'b00011111000: dataA <= 32'b10011011101110000010010110101110;
11'b00011111001: dataA <= 32'b00001001010000011111010011011001;
11'b00011111010: dataA <= 32'b01011111000010001111101010010011;
11'b00011111011: dataA <= 32'b00000011101100001100011010011011;
11'b00011111100: dataA <= 32'b00010111010001101110011010101011;
11'b00011111101: dataA <= 32'b00001100010111110101000001110100;
11'b00011111110: dataA <= 32'b10001010100010110011100111110110;
11'b00011111111: dataA <= 32'b00001111001111110000110001010001;
11'b00100000000: dataA <= 32'b11100111101011110101001011110001;
11'b00100000001: dataA <= 32'b00001101111001101011001110111101;
11'b00100000010: dataA <= 32'b10101000111011001011001011110100;
11'b00100000011: dataA <= 32'b00000100001100001100010110011111;
11'b00100000100: dataA <= 32'b01000111100001101100110110011001;
11'b00100000101: dataA <= 32'b00000000110101000101000000011101;
11'b00100000110: dataA <= 32'b11010111010011110011011100001010;
11'b00100000111: dataA <= 32'b00000000110000000110101101101011;
11'b00100001000: dataA <= 32'b01101111110101010101110011111011;
11'b00100001001: dataA <= 32'b00001010101111101010100111011110;
11'b00100001010: dataA <= 32'b00010000001001101110011000000100;
11'b00100001011: dataA <= 32'b00000101010001010010101101010001;
11'b00100001100: dataA <= 32'b01100001000010110100101001110110;
11'b00100001101: dataA <= 32'b00001011111101110100011010010101;
11'b00100001110: dataA <= 32'b00101100010100111110000011110011;
11'b00100001111: dataA <= 32'b00000111011100011101011111010001;
11'b00100010000: dataA <= 32'b01100010011111011010111100100100;
11'b00100010001: dataA <= 32'b00001100011011101011011010001011;
11'b00100010010: dataA <= 32'b11001010010111101101101100011010;
11'b00100010011: dataA <= 32'b00000011110010000110110100110110;
11'b00100010100: dataA <= 32'b10100011010010110010111000011010;
11'b00100010101: dataA <= 32'b00000010001000000110110110000110;
11'b00100010110: dataA <= 32'b00001100111111110010111001111010;
11'b00100010111: dataA <= 32'b00001001000001011011010000111101;
11'b00100011000: dataA <= 32'b11100110011101101101100110010001;
11'b00100011001: dataA <= 32'b00000100011011001001100110010110;
11'b00100011010: dataA <= 32'b10000101010101000010000011010100;
11'b00100011011: dataA <= 32'b00001110110101110100111100111100;
11'b00100011100: dataA <= 32'b10010100100011110100001011010010;
11'b00100011101: dataA <= 32'b00000001001000001100010001011011;
11'b00100011110: dataA <= 32'b00100001011011100001111000010011;
11'b00100011111: dataA <= 32'b00000101111100011000110010010100;
11'b00100100000: dataA <= 32'b00011011100011110011011100110000;
11'b00100100001: dataA <= 32'b00000011101001000111100001111011;
11'b00100100010: dataA <= 32'b01011111111010111001111001011101;
11'b00100100011: dataA <= 32'b00001001010110101000100010010011;
11'b00100100100: dataA <= 32'b00100110000101010101010100100010;
11'b00100100101: dataA <= 32'b00001011010101101001100110000110;
11'b00100100110: dataA <= 32'b10001001001011001011101100001001;
11'b00100100111: dataA <= 32'b00000110100101010000001101001100;
11'b00100101000: dataA <= 32'b11010100001010011110111001010110;
11'b00100101001: dataA <= 32'b00001011101010100111001001001001;
11'b00100101010: dataA <= 32'b00010001101100110101100010111010;
11'b00100101011: dataA <= 32'b00001010111101101101100101010100;
11'b00100101100: dataA <= 32'b11110011100001110100110111001110;
11'b00100101101: dataA <= 32'b00000101001010000011010111010110;
11'b00100101110: dataA <= 32'b01100010100101000110110101000001;
11'b00100101111: dataA <= 32'b00001001001001011110110110100000;
11'b00100110000: dataA <= 32'b01010101011001100100100110000110;
11'b00100110001: dataA <= 32'b00001011110001101100110001010111;
11'b00100110010: dataA <= 32'b01011011000110111101011010001111;
11'b00100110011: dataA <= 32'b00001110000111011111111001111111;
11'b00100110100: dataA <= 32'b11101110110001111011100101011100;
11'b00100110101: dataA <= 32'b00001001110111100111001011010110;
11'b00100110110: dataA <= 32'b10010100001101001011010100010010;
11'b00100110111: dataA <= 32'b00000000110100001000011100111101;
11'b00100111000: dataA <= 32'b00011111111010111110011011110100;
11'b00100111001: dataA <= 32'b00000011001011001000111110011010;
11'b00100111010: dataA <= 32'b11011011011110001000010101111100;
11'b00100111011: dataA <= 32'b00000000110001000101011110001001;
11'b00100111100: dataA <= 32'b01011010100101100011110010111010;
11'b00100111101: dataA <= 32'b00000110010110011110000101011110;
11'b00100111110: dataA <= 32'b00101011011011110011011110000111;
11'b00100111111: dataA <= 32'b00001000101001100010000111110101;
11'b00101000000: dataA <= 32'b11010010100101000101100100010000;
11'b00101000001: dataA <= 32'b00000110101010010101000001000101;
11'b00101000010: dataA <= 32'b10100111100011001100101101000100;
11'b00101000011: dataA <= 32'b00000111011100100010010111000110;
11'b00101000100: dataA <= 32'b10011111110111000101111010111100;
11'b00101000101: dataA <= 32'b00001101111010101001111010001101;
11'b00101000110: dataA <= 32'b10011000110110101111101010100010;
11'b00101000111: dataA <= 32'b00001010111101100101110101100100;
11'b00101001000: dataA <= 32'b00100110111001010011010000101100;
11'b00101001001: dataA <= 32'b00000011100101001001011110010110;
11'b00101001010: dataA <= 32'b10101110100111001110011101001100;
11'b00101001011: dataA <= 32'b00000101101001010110010010100111;
11'b00101001100: dataA <= 32'b11101000111001000010110011110000;
11'b00101001101: dataA <= 32'b00001010100101100001010111100001;
11'b00101001110: dataA <= 32'b10100011101101110010010110101111;
11'b00101001111: dataA <= 32'b00001001001111100011010010110000;
11'b00101010000: dataA <= 32'b00011111000010111111011010110001;
11'b00101010001: dataA <= 32'b00000011010000000110101010001011;
11'b00101010010: dataA <= 32'b00011011010110001110011001101001;
11'b00101010011: dataA <= 32'b00001101010100110010110001110100;
11'b00101010100: dataA <= 32'b01000110110110100010111000110110;
11'b00101010101: dataA <= 32'b00001110101001101100100100111010;
11'b00101010110: dataA <= 32'b11101111100011110011111011101110;
11'b00101010111: dataA <= 32'b00001111010100101101000111001100;
11'b00101011000: dataA <= 32'b00011100101101100001101010001000;
11'b00101011001: dataA <= 32'b00000110010111001011100111110011;
11'b00101011010: dataA <= 32'b00110001110010011100101100110011;
11'b00101011011: dataA <= 32'b00001010111110100001110110101111;
11'b00101011100: dataA <= 32'b10101001010001101000010101000111;
11'b00101011101: dataA <= 32'b00001000011110010111110001111100;
11'b00101011110: dataA <= 32'b00111010100010111101011101111000;
11'b00101011111: dataA <= 32'b00000111101010010010101011001001;
11'b00101100000: dataA <= 32'b01000101011111001100100010001111;
11'b00101100001: dataA <= 32'b00001000110101010111011000100101;
11'b00101100010: dataA <= 32'b01100000111110010010011011001100;
11'b00101100011: dataA <= 32'b00001110101000001100010110101011;
11'b00101100100: dataA <= 32'b01001010100111000110001001111000;
11'b00101100101: dataA <= 32'b00001110010001101111000100100001;
11'b00101100110: dataA <= 32'b10001110111001011001000010000110;
11'b00101100111: dataA <= 32'b00001101100111101100101001101011;
11'b00101101000: dataA <= 32'b01001011101010110000101101000111;
11'b00101101001: dataA <= 32'b00001001011000011011110011011110;
11'b00101101010: dataA <= 32'b11101000111001011010011101001111;
11'b00101101011: dataA <= 32'b00000100011011011011110011010011;
11'b00101101100: dataA <= 32'b00011111100101011000011101001100;
11'b00101101101: dataA <= 32'b00000000101101101001001010100110;
11'b00101101110: dataA <= 32'b01001110110010110100101000110011;
11'b00101101111: dataA <= 32'b00001101110111110011101111011011;
11'b00101110000: dataA <= 32'b00101011110101000101111010011001;
11'b00101110001: dataA <= 32'b00001010100010011110010110010110;
11'b00101110010: dataA <= 32'b00010001010110000000011001001001;
11'b00101110011: dataA <= 32'b00000100011101001001100101110101;
11'b00101110100: dataA <= 32'b01101100111100111000111001101111;
11'b00101110101: dataA <= 32'b00001110010100011001001110000011;
11'b00101110110: dataA <= 32'b00110001001001101000011000000110;
11'b00101110111: dataA <= 32'b00000100111000110001110001100100;
11'b00101111000: dataA <= 32'b01111101000000111010001110101101;
11'b00101111001: dataA <= 32'b00001011001101010000101101101011;
11'b00101111010: dataA <= 32'b11000010110010101101010001010110;
11'b00101111011: dataA <= 32'b00001010101001110010101111000011;
11'b00101111100: dataA <= 32'b10100101101101110001100100100111;
11'b00101111101: dataA <= 32'b00000010110010000111011110010101;
11'b00101111110: dataA <= 32'b10000101010111011011001011001101;
11'b00101111111: dataA <= 32'b00000101001000100100110000111101;
11'b00110000000: dataA <= 32'b01110111011110110110011101011010;
11'b00110000001: dataA <= 32'b00001110101010110010100110000101;
11'b00110000010: dataA <= 32'b01110000011010011100010111010001;
11'b00110000011: dataA <= 32'b00000101010101101011111011011001;
11'b00110000100: dataA <= 32'b11010010111011011101110000110101;
11'b00110000101: dataA <= 32'b00000100101101011011000000001010;
11'b00110000110: dataA <= 32'b01101101010110010100110011010011;
11'b00110000111: dataA <= 32'b00001000101000011000100111101101;
11'b00110001000: dataA <= 32'b00100011001010101010000111101011;
11'b00110001001: dataA <= 32'b00000011100011111101000011101100;
11'b00110001010: dataA <= 32'b01011000100001110100001110010101;
11'b00110001011: dataA <= 32'b00001011101100100100110011011001;
11'b00110001100: dataA <= 32'b00000111010101101101101001010111;
11'b00110001101: dataA <= 32'b00001010011110001111101110110110;
11'b00110001110: dataA <= 32'b00111101000011001010001010001000;
11'b00110001111: dataA <= 32'b00000101111001011111101101000011;
11'b00110010000: dataA <= 32'b10101111001000001011101110010100;
11'b00110010001: dataA <= 32'b00001000111110101111110100111011;
11'b00110010010: dataA <= 32'b00010011001001111100111101011010;
11'b00110010011: dataA <= 32'b00001011010011000011000011001101;
11'b00110010100: dataA <= 32'b01101100101001101000010011100011;
11'b00110010101: dataA <= 32'b00000100101110000010111010100000;
11'b00110010110: dataA <= 32'b11010011011010110101111000010111;
11'b00110010111: dataA <= 32'b00000101010010100001010110111101;
11'b00110011000: dataA <= 32'b11110000110010010001100010000101;
11'b00110011001: dataA <= 32'b00001110010001001010111011010001;
11'b00110011010: dataA <= 32'b10111011000010111001111110001010;
11'b00110011011: dataA <= 32'b00001101000100111100101110110011;
11'b00110011100: dataA <= 32'b11011011001111110010100001001010;
11'b00110011101: dataA <= 32'b00001110101010111010110110010100;
11'b00110011110: dataA <= 32'b01011100110001101101010110011110;
11'b00110011111: dataA <= 32'b00000010111000101111101111000011;
11'b00110100000: dataA <= 32'b11010010100011001001100110000101;
11'b00110100001: dataA <= 32'b00000100110100001001010011110010;
11'b00110100010: dataA <= 32'b11011100101101011101111000011000;
11'b00110100011: dataA <= 32'b00000010101010101010111100111000;
11'b00110100100: dataA <= 32'b01110110111001001100010111110010;
11'b00110100101: dataA <= 32'b00000111101101101000111000010010;
11'b00110100110: dataA <= 32'b10100001000011101010001000101010;
11'b00110100111: dataA <= 32'b00001000011001010101110001100011;
11'b00110101000: dataA <= 32'b01101011001011001011100100101100;
11'b00110101001: dataA <= 32'b00001010000101011000011010000100;
11'b00110101010: dataA <= 32'b00011011110001011010111011001110;
11'b00110101011: dataA <= 32'b00000100100010010010100101001110;
11'b00110101100: dataA <= 32'b10110000100001111000010111001000;
11'b00110101101: dataA <= 32'b00001010000001100010100110011001;
11'b00110101110: dataA <= 32'b10100000101110000001011011001011;
11'b00110101111: dataA <= 32'b00000100110101000101010011110100;
11'b00110110000: dataA <= 32'b01100101111010010100111011110111;
11'b00110110001: dataA <= 32'b00000111111110010111110010000111;
11'b00110110010: dataA <= 32'b10100011011010011000010111000110;
11'b00110110011: dataA <= 32'b00000101011101001111100101110100;
11'b00110110100: dataA <= 32'b00111100111010100101111011111100;
11'b00110110101: dataA <= 32'b00001000101011011000100011101010;
11'b00110110110: dataA <= 32'b01000011000110111101100010101011;
11'b00110110111: dataA <= 32'b00000111110101010011010000011100;
11'b00110111000: dataA <= 32'b11100000111110100010101011101111;
11'b00110111001: dataA <= 32'b00001111001110010110001010110011;
11'b00110111010: dataA <= 32'b10010010011010100110110111111001;
11'b00110111011: dataA <= 32'b00001101110110101101010001001000;
11'b00110111100: dataA <= 32'b01010000101001111000110100000010;
11'b00110111101: dataA <= 32'b00001111001100110000110001110011;
11'b00110111110: dataA <= 32'b01000101011011011001101110101100;
11'b00110111111: dataA <= 32'b00000111011000010001101010111111;
11'b00111000000: dataA <= 32'b11101001000001101010001100110011;
11'b00111000001: dataA <= 32'b00000010011000010001101011001100;
11'b00111000010: dataA <= 32'b01010111100010001000011101110000;
11'b00111000011: dataA <= 32'b00000001100111100111010010001110;
11'b00111000100: dataA <= 32'b01010010100110101101000111110011;
11'b00111000101: dataA <= 32'b00001100011011101001111011011100;
11'b00111000110: dataA <= 32'b00011111111000110101000111111010;
11'b00111000111: dataA <= 32'b00001101000101100110011001110110;
11'b00111001000: dataA <= 32'b11001111001010110000101010001010;
11'b00111001001: dataA <= 32'b00000010011001000011010001100100;
11'b00111001010: dataA <= 32'b01101101000101101000011001110000;
11'b00111001011: dataA <= 32'b00001100111000010111000110001011;
11'b00111001100: dataA <= 32'b11101101010110011000011010000111;
11'b00111001101: dataA <= 32'b00000011010101100101111001100011;
11'b00111001110: dataA <= 32'b00111011011001011001011110110011;
11'b00111001111: dataA <= 32'b00001011110000010110100101110011;
11'b00111010000: dataA <= 32'b10001000011010010101100000110000;
11'b00111010001: dataA <= 32'b00001011101100110101000010111100;
11'b00111010010: dataA <= 32'b11011101101110010001100110100101;
11'b00111010011: dataA <= 32'b00000010001110000011001001111101;
11'b00111010100: dataA <= 32'b10000010111111100100011011110000;
11'b00111010101: dataA <= 32'b00000110100111100110110100101100;
11'b00111010110: dataA <= 32'b01110001101110010110111010111101;
11'b00111010111: dataA <= 32'b00001111001111110110110101110101;
11'b00111011000: dataA <= 32'b10110110101010010100110111010001;
11'b00111011001: dataA <= 32'b00000100110010011111111011110010;
11'b00111011010: dataA <= 32'b10010100110011000110110000101111;
11'b00111011011: dataA <= 32'b00000101001011011010111100100001;
11'b00111011100: dataA <= 32'b10100111011110000101000010101111;
11'b00111011101: dataA <= 32'b00001010001001011110100011010110;
11'b00111011110: dataA <= 32'b01100001001010111010111000101100;
11'b00111011111: dataA <= 32'b00000110100001111011011011011101;
11'b00111100000: dataA <= 32'b10011110011101110100001100111001;
11'b00111100001: dataA <= 32'b00001100001111100110110111110010;
11'b00111100010: dataA <= 32'b10000101000001011101010111111000;
11'b00111100011: dataA <= 32'b00000111011110000111011110010110;
11'b00111100100: dataA <= 32'b01111011011011011011001011001011;
11'b00111100101: dataA <= 32'b00000011110110010111101001010010;
11'b00111100110: dataA <= 32'b10101101010100011010001100111000;
11'b00111100111: dataA <= 32'b00000110011110100011111001000010;
11'b00111101000: dataA <= 32'b00010000111101101100111010111101;
11'b00111101001: dataA <= 32'b00001010010101000010101110110110;
11'b00111101010: dataA <= 32'b00110000110010011000010110100001;
11'b00111101011: dataA <= 32'b00000101001100000110100011001001;
11'b00111101100: dataA <= 32'b01001111001110011110010110110110;
11'b00111101101: dataA <= 32'b00000100110000011101010010100110;
11'b00111101110: dataA <= 32'b00110011000010110010000100100010;
11'b00111101111: dataA <= 32'b00001101110110001100101011101011;
11'b00111110000: dataA <= 32'b00110111010111010010111110101111;
11'b00111110001: dataA <= 32'b00001110101001111101000110110100;
11'b00111110010: dataA <= 32'b00011001001011110100000010100101;
11'b00111110011: dataA <= 32'b00001111010000111011001110000101;
11'b00111110100: dataA <= 32'b01100000110001011101000011011011;
11'b00111110101: dataA <= 32'b00000001010011100101110111000100;
11'b00111110110: dataA <= 32'b01011000011011100010111000000100;
11'b00111110111: dataA <= 32'b00000100010010000111000011110100;
11'b00111111000: dataA <= 32'b01100000101101001101000110110111;
11'b00111111001: dataA <= 32'b00000100000111101011000101101000;
11'b00111111010: dataA <= 32'b00110111001001001011110111010010;
11'b00111111011: dataA <= 32'b00001000001101101001000000110001;
11'b00111111100: dataA <= 32'b00100001000011110011101001101011;
11'b00111111101: dataA <= 32'b00000110011000001101100101101011;
11'b00111111110: dataA <= 32'b01101001010011001100100101101010;
11'b00111111111: dataA <= 32'b00001011100111100000010110000100;
11'b01000000000: dataA <= 32'b01010001101001110010011011010000;
11'b01000000001: dataA <= 32'b00000111100001011000011100110101;
11'b01000000010: dataA <= 32'b00110100110010100000011000101000;
11'b01000000011: dataA <= 32'b00001100100100100110101010111010;
11'b01000000100: dataA <= 32'b11100100110010100001101100001110;
11'b01000000101: dataA <= 32'b00000100010010000010111011100101;
11'b01000000110: dataA <= 32'b00011011111010000101001001111001;
11'b01000000111: dataA <= 32'b00000100111101001101100101011111;
11'b01000001000: dataA <= 32'b01011111011011000000111000100110;
11'b01000001001: dataA <= 32'b00000010111010001001010101101100;
11'b01000001010: dataA <= 32'b10111101010010001110001001011110;
11'b01000001011: dataA <= 32'b00001001101100011110011111110011;
11'b01000001100: dataA <= 32'b00000010110010100110000100000111;
11'b01000001101: dataA <= 32'b00000110110101010001000100011011;
11'b01000001110: dataA <= 32'b01100000111110110011001011110010;
11'b01000001111: dataA <= 32'b00001111010100100010000110110100;
11'b01000010000: dataA <= 32'b01011010010001111111000110011000;
11'b01000010001: dataA <= 32'b00001100011010101001011001111000;
11'b01000010010: dataA <= 32'b00010100100010100001000111000001;
11'b01000010011: dataA <= 32'b00001111010010110001000001111011;
11'b01000010100: dataA <= 32'b10000011000011110010111110110001;
11'b01000010101: dataA <= 32'b00000101110111001011011110001111;
11'b01000010110: dataA <= 32'b10100111001010000010001100010110;
11'b01000010111: dataA <= 32'b00000001010011001011011111000101;
11'b01000011000: dataA <= 32'b00010011010110111000101101010100;
11'b01000011001: dataA <= 32'b00000011100011100011010101101110;
11'b01000011010: dataA <= 32'b10011000011110011101100111010011;
11'b01000011011: dataA <= 32'b00001001111101011101111011010101;
11'b01000011100: dataA <= 32'b11010101110100101100000101111001;
11'b01000011101: dataA <= 32'b00001110101010101110100001011101;
11'b01000011110: dataA <= 32'b01001100111011011001101011001100;
11'b01000011111: dataA <= 32'b00000000110011000010111001011100;
11'b01000100000: dataA <= 32'b10101001001110010000011001010001;
11'b01000100001: dataA <= 32'b00001010111011010110111110010011;
11'b01000100010: dataA <= 32'b10101001100011000000111011001010;
11'b01000100011: dataA <= 32'b00000010010001011011111001101011;
11'b01000100100: dataA <= 32'b00110011101101111001001101111000;
11'b01000100101: dataA <= 32'b00001011010010011100011101111011;
11'b01000100110: dataA <= 32'b01010000001110000101110000101010;
11'b01000100111: dataA <= 32'b00001100001111110011010010110101;
11'b01000101000: dataA <= 32'b10010011101010101010001000100101;
11'b01000101001: dataA <= 32'b00000011001010000010110001101101;
11'b01000101010: dataA <= 32'b10000100101011011101011011010010;
11'b01000101011: dataA <= 32'b00001000100110101000111100101011;
11'b01000101100: dataA <= 32'b00100111110101101110110111111110;
11'b01000101101: dataA <= 32'b00001110110101110111001001100101;
11'b01000101110: dataA <= 32'b00111000111010001100110110110000;
11'b01000101111: dataA <= 32'b00000100010000010011110111110100;
11'b01000110000: dataA <= 32'b10011000101010011111010001001001;
11'b01000110001: dataA <= 32'b00000110001001011100111001001000;
11'b01000110010: dataA <= 32'b01100001100001111101000011001011;
11'b01000110011: dataA <= 32'b00001011001011100100100010101111;
11'b01000110100: dataA <= 32'b01011111001011000011101001001100;
11'b01000110101: dataA <= 32'b00001001000001110011101111000110;
11'b01000110110: dataA <= 32'b00100110011101110011111010011100;
11'b01000110111: dataA <= 32'b00001100010011101000111111110100;
11'b01000111000: dataA <= 32'b10000110101101001100110110010111;
11'b01000111001: dataA <= 32'b00000100011101000011001001110110;
11'b01000111010: dataA <= 32'b00110011101111011100011100001110;
11'b01000111011: dataA <= 32'b00000011010011001111011101101010;
11'b01000111100: dataA <= 32'b00100111011100110001001010111011;
11'b01000111101: dataA <= 32'b00000011011011010111111001010010;
11'b01000111110: dataA <= 32'b01010010110101100100100111111110;
11'b01000111111: dataA <= 32'b00001001010110001000011010011110;
11'b01001000000: dataA <= 32'b01110001000011000000111001000001;
11'b01001000001: dataA <= 32'b00000110001010001100010011101010;
11'b01001000010: dataA <= 32'b10001101000001111110010101110101;
11'b01001000011: dataA <= 32'b00000100101110011001001110000110;
11'b01001000100: dataA <= 32'b01110001001111000010110111100001;
11'b01001000101: dataA <= 32'b00001100011010010010011111101100;
11'b01001000110: dataA <= 32'b11110001100111011011111110010100;
11'b01001000111: dataA <= 32'b00001111001111111011011010101100;
11'b01001001000: dataA <= 32'b00010111000011101101100101000010;
11'b01001001001: dataA <= 32'b00001110110101110111100001111101;
11'b01001001010: dataA <= 32'b00100010110001010100100001110111;
11'b01001001011: dataA <= 32'b00000001001110011011110110111101;
11'b01001001100: dataA <= 32'b11100000011011101100001010000101;
11'b01001001101: dataA <= 32'b00000100001111001000101111101101;
11'b01001001110: dataA <= 32'b01100100110000111100010101010110;
11'b01001001111: dataA <= 32'b00000110000101101001001110010000;
11'b01001010000: dataA <= 32'b01110011011001010011000110110001;
11'b01001010001: dataA <= 32'b00001000101110100111001001011000;
11'b01001010010: dataA <= 32'b00100001000011110101001010001100;
11'b01001010011: dataA <= 32'b00000100110110000111010001110011;
11'b01001010100: dataA <= 32'b01100101010110111101010110101001;
11'b01001010101: dataA <= 32'b00001101001011101000011001111100;
11'b01001010110: dataA <= 32'b01001011011110000010011010110011;
11'b01001010111: dataA <= 32'b00001010100001011110011000100100;
11'b01001011000: dataA <= 32'b00110111000011001001001010001001;
11'b01001011001: dataA <= 32'b00001110101001101010110011001011;
11'b01001011010: dataA <= 32'b00100110110110111010011100010001;
11'b01001011011: dataA <= 32'b00000011101111000110100111000111;
11'b01001011100: dataA <= 32'b01001111110001110101000111111010;
11'b01001011101: dataA <= 32'b00000010011010000111010100110110;
11'b01001011110: dataA <= 32'b00011011010111100001111010100111;
11'b01001011111: dataA <= 32'b00000001010101000101000001101100;
11'b01001100000: dataA <= 32'b00110111100101101110000110011101;
11'b01001100001: dataA <= 32'b00001010001110100100100011110101;
11'b01001100010: dataA <= 32'b11001000011010000110100101100101;
11'b01001100011: dataA <= 32'b00000101110011010000111000110001;
11'b01001100100: dataA <= 32'b00100000111110111011111011010100;
11'b01001100101: dataA <= 32'b00001101111001101100001110100101;
11'b01001100110: dataA <= 32'b01100010010001011110110100110110;
11'b01001100111: dataA <= 32'b00001001111100100011011110101000;
11'b01001101000: dataA <= 32'b00011100011111000001111010000001;
11'b01001101001: dataA <= 32'b00001110010111101111001110000011;
11'b01001101010: dataA <= 32'b10000010101011110100001101110110;
11'b01001101011: dataA <= 32'b00000100010101000111001001011111;
11'b01001101100: dataA <= 32'b01100101001110011010011010011001;
11'b01001101101: dataA <= 32'b00000001001101000111001010100110;
11'b01001101110: dataA <= 32'b11001111001011011001101011111000;
11'b01001101111: dataA <= 32'b00000110100001011111010101010101;
11'b01001110000: dataA <= 32'b01100000011010000101110110110010;
11'b01001110001: dataA <= 32'b00000110111101010001110110111110;
11'b01001110010: dataA <= 32'b01001011101000110010110100010111;
11'b01001110011: dataA <= 32'b00001111010000110010110001000101;
11'b01001110100: dataA <= 32'b11001110101111110010111011101111;
11'b01001110101: dataA <= 32'b00000000101110000100100001010011;
11'b01001110110: dataA <= 32'b11100111010111000000111000110010;
11'b01001110111: dataA <= 32'b00001000011101010110110110010011;
11'b01001111000: dataA <= 32'b01100001100111100001111100001101;
11'b01001111001: dataA <= 32'b00000010101101001111110001110011;
11'b01001111010: dataA <= 32'b00101001111010011001011011111011;
11'b01001111011: dataA <= 32'b00001010110101100010011110001011;
11'b01001111100: dataA <= 32'b11011100000101101101100010000101;
11'b01001111101: dataA <= 32'b00001011110010101111011110011101;
11'b01001111110: dataA <= 32'b01001101011111000010111010100110;
11'b01001111111: dataA <= 32'b00000100100111001000011101010101;
11'b01010000000: dataA <= 32'b10001010010111000110011010110101;
11'b01010000001: dataA <= 32'b00001010000111101001000100110010;
11'b01010000010: dataA <= 32'b10011011110101001110010101011101;
11'b01010000011: dataA <= 32'b00001101011010110011011001011100;
11'b01010000100: dataA <= 32'b10110111001101111101000110101111;
11'b01010000101: dataA <= 32'b00000100101101001001101011101101;
11'b01010000110: dataA <= 32'b01011100100101101111010010100100;
11'b01010000111: dataA <= 32'b00000111101000011100111001111000;
11'b01010001000: dataA <= 32'b10011011011101101100110100101000;
11'b01010001001: dataA <= 32'b00001011101110101000100101111111;
11'b01010001010: dataA <= 32'b00011101001011000100101001101110;
11'b01010001011: dataA <= 32'b00001100000011101001111010100111;
11'b01010001100: dataA <= 32'b10101010100101110011110111111101;
11'b01010001101: dataA <= 32'b00001011010101101001000111101101;
11'b01010001110: dataA <= 32'b01001100011001000100000100110101;
11'b01010001111: dataA <= 32'b00000010011001000100110001010110;
11'b01010010000: dataA <= 32'b11101001111011010101101100010001;
11'b01010010001: dataA <= 32'b00000010101111001011010010000001;
11'b01010010010: dataA <= 32'b11100001100001100000011000011101;
11'b01010010011: dataA <= 32'b00000001010111001101101101110001;
11'b01010010100: dataA <= 32'b10010100101001100100000101011101;
11'b01010010101: dataA <= 32'b00000111110111010010001001111110;
11'b01010010110: dataA <= 32'b11101111001111100001111100000011;
11'b01010010111: dataA <= 32'b00000111001001011000000111110011;
11'b01010011000: dataA <= 32'b01001110110001011110010100110011;
11'b01010011001: dataA <= 32'b00000101101011010111000101011110;
11'b01010011010: dataA <= 32'b10101101011011010011111010100001;
11'b01010011011: dataA <= 32'b00001001111100011000010111011101;
11'b01010011100: dataA <= 32'b01101001110011010100111100111001;
11'b01010011101: dataA <= 32'b00001111010101110011101110100101;
11'b01010011110: dataA <= 32'b11010110111011010110101000000001;
11'b01010011111: dataA <= 32'b00001101011010101111101101101100;
11'b01010100000: dataA <= 32'b11100100110101001100000000110001;
11'b01010100001: dataA <= 32'b00000010001001010001101110101101;
11'b01010100010: dataA <= 32'b11101000011011100101011100001000;
11'b01010100011: dataA <= 32'b00000100101100001110011111001110;
11'b01010100100: dataA <= 32'b11100110110100111011100100010011;
11'b01010100101: dataA <= 32'b00001000000100100101010011000000;
11'b01010100110: dataA <= 32'b01101101101001011010100110110000;
11'b01010100111: dataA <= 32'b00001000101110100101001110000000;
11'b01010101000: dataA <= 32'b11100001000011011110011010101110;
11'b01010101001: dataA <= 32'b00000011110011000100111110000010;
11'b01010101010: dataA <= 32'b01100001011010100110001000001000;
11'b01010101011: dataA <= 32'b00001101101111101110100101111100;
11'b01010101100: dataA <= 32'b01000111001010010010101010010101;
11'b01010101101: dataA <= 32'b00001101000100100110011100101011;
11'b01010101110: dataA <= 32'b00110101010111101010011011001011;
11'b01010101111: dataA <= 32'b00001111001111101100111011010100;
11'b01010110000: dataA <= 32'b11011010110001001010001000100111;
11'b01010110001: dataA <= 32'b00000111111000010011110011100001;
11'b01010110010: dataA <= 32'b01111001100010100100011101010000;
11'b01010110011: dataA <= 32'b00001101011011101011110011001110;
11'b01010110100: dataA <= 32'b10101011001000111000110011101010;
11'b01010110101: dataA <= 32'b00001010111101100001110110000100;
11'b01010110110: dataA <= 32'b01110010010011000100101110110011;
11'b01010110111: dataA <= 32'b00000111001011010000110110100000;
11'b01010111000: dataA <= 32'b01001101101111010011110010110100;
11'b01010111001: dataA <= 32'b00001001110100011101011100111110;
11'b01010111010: dataA <= 32'b11011110111101111010001010001001;
11'b01010111011: dataA <= 32'b00001100100100000110100110100010;
11'b01010111100: dataA <= 32'b10001000111011011101001011010110;
11'b01010111101: dataA <= 32'b00001110001100101110111000001010;
11'b01010111110: dataA <= 32'b11001111000100111001110000101011;
11'b01010111111: dataA <= 32'b00001011100011100110100001100011;
11'b01011000000: dataA <= 32'b00010101111010000000011011000100;
11'b01011000001: dataA <= 32'b00001010110111100101110011110101;
11'b01011000010: dataA <= 32'b11100110110101001011001100101011;
11'b01011000011: dataA <= 32'b00000110111101100101110011001010;
11'b01011000100: dataA <= 32'b01100101100000110001001100001000;
11'b01011000101: dataA <= 32'b00000000110010101011000010111101;
11'b01011000110: dataA <= 32'b00001100111110111011111001010010;
11'b01011000111: dataA <= 32'b00001110110010111011011111001010;
11'b01011001000: dataA <= 32'b11110101101001011110011011110111;
11'b01011001001: dataA <= 32'b00001000000001011000011010101101;
11'b01011001010: dataA <= 32'b01010111100001011000010111101000;
11'b01011001011: dataA <= 32'b00000111011110010001110101111101;
11'b01011001100: dataA <= 32'b01101010110000011001111001001110;
11'b01011001101: dataA <= 32'b00001110101111011011010001111011;
11'b01011001110: dataA <= 32'b01110010111100111000110110100111;
11'b01011001111: dataA <= 32'b00000110111010111001100001101100;
11'b01011010000: dataA <= 32'b10111100101100101011001101101000;
11'b01011010001: dataA <= 32'b00001010101010001110111001100011;
11'b01011010010: dataA <= 32'b00000011000110110100100010111011;
11'b01011010011: dataA <= 32'b00001001001000101110100010111011;
11'b01011010100: dataA <= 32'b01101111100101011001110011001010;
11'b01011010101: dataA <= 32'b00000011110110001111101110101101;
11'b01011010110: dataA <= 32'b01001011101011001001111010101010;
11'b01011010111: dataA <= 32'b00000011101011100010101101010110;
11'b01011011000: dataA <= 32'b00111011001011001101101110110101;
11'b01011011001: dataA <= 32'b00001101000101101100011010010101;
11'b01011011010: dataA <= 32'b10100110010010100100000111110010;
11'b01011011011: dataA <= 32'b00000110110110110101101110110000;
11'b01011011100: dataA <= 32'b00010011000111101100100010011010;
11'b01011011101: dataA <= 32'b00000100010000011101000100001100;
11'b01011011110: dataA <= 32'b00101111001010011100100100010110;
11'b01011011111: dataA <= 32'b00000111001000010010101111110100;
11'b01011100000: dataA <= 32'b11100101000110010001110111001100;
11'b01011100001: dataA <= 32'b00000001100111111100101111100010;
11'b01011100010: dataA <= 32'b10010010101001111100011110110000;
11'b01011100011: dataA <= 32'b00001010101001100010101110110000;
11'b01011100100: dataA <= 32'b01001101100110000101111010110110;
11'b01011100101: dataA <= 32'b00001100111011011001110111001101;
11'b01011100110: dataA <= 32'b11111100101110110001011000100111;
11'b01011100111: dataA <= 32'b00000111111010101001101000111011;
11'b01011101000: dataA <= 32'b01110000111100001100111110101111;
11'b01011101001: dataA <= 32'b00001011111101110111100100111100;
11'b01011101010: dataA <= 32'b00010101010110000100111110110101;
11'b01011101011: dataA <= 32'b00001011110000000101011011010100;
11'b01011101100: dataA <= 32'b01100110100000111000110001100111;
11'b01011101101: dataA <= 32'b00000100110001000011001101111000;
11'b01011101110: dataA <= 32'b00011001100011001101001001110110;
11'b01011101111: dataA <= 32'b00000101110100100011010011001101;
11'b01011110000: dataA <= 32'b00101100100101111001010000101010;
11'b01011110001: dataA <= 32'b00001110001100001011001110110001;
11'b01011110010: dataA <= 32'b11111000101110011001011100100110;
11'b01011110011: dataA <= 32'b00001010100001110110011010101010;
11'b01011110100: dataA <= 32'b10011101010011010001010000101111;
11'b01011110101: dataA <= 32'b00001101000101110110100010011100;
11'b01011110110: dataA <= 32'b10011010110110000101101000111110;
11'b01011110111: dataA <= 32'b00000100111011110111011110111010;
11'b01011111000: dataA <= 32'b10001100101110101000110100000111;
11'b01011111001: dataA <= 32'b00000110010110001111100011011001;
11'b01011111010: dataA <= 32'b11011010110001110110001001110111;
11'b01011111011: dataA <= 32'b00000010001111101000110100011001;
11'b01011111100: dataA <= 32'b11110100100101010101001000010010;
11'b01011111101: dataA <= 32'b00000111001110100110110100001011;
11'b01011111110: dataA <= 32'b11100000111111001001000111001010;
11'b01011111111: dataA <= 32'b00001001111000011111110101011011;
11'b01100000000: dataA <= 32'b00101100111111000010110100001111;
11'b01100000001: dataA <= 32'b00000111100100010010100010001100;
11'b01100000010: dataA <= 32'b10100101110001010011011010101011;
11'b01100000011: dataA <= 32'b00000010000101001110110001101110;
11'b01100000100: dataA <= 32'b01101010010101001000100101101001;
11'b01100000101: dataA <= 32'b00000111100001011100100110000001;
11'b01100000110: dataA <= 32'b11011000110100110010110111000111;
11'b01100000111: dataA <= 32'b00001001010111011101111010111000;
11'b01100001000: dataA <= 32'b00111101001010100011111100101100;
11'b01100001001: dataA <= 32'b00001110110110110011100111100101;
11'b01100001010: dataA <= 32'b10101101000000011001110011001110;
11'b01100001011: dataA <= 32'b00001101011010101011101110001100;
11'b01100001100: dataA <= 32'b01101000000111000011101111001101;
11'b01100001101: dataA <= 32'b00000110001100001111000001110000;
11'b01100001110: dataA <= 32'b00011001111011000010110011110111;
11'b01100001111: dataA <= 32'b00001010110010100011011101100111;
11'b01100010000: dataA <= 32'b01011110111101100010011001001000;
11'b01100010001: dataA <= 32'b00001010000001000010111010001010;
11'b01100010010: dataA <= 32'b00001001001011100100001100010011;
11'b01100010011: dataA <= 32'b00001101000111101100101100001100;
11'b01100010100: dataA <= 32'b00010001010100100010110000110001;
11'b01100010101: dataA <= 32'b00001001000001100000011101100100;
11'b01100010110: dataA <= 32'b10100001111001011000011000100010;
11'b01100010111: dataA <= 32'b00001011110100101111101011110011;
11'b01100011000: dataA <= 32'b11100100110001000011111011000111;
11'b01100011001: dataA <= 32'b00001001111101101111101010110001;
11'b01100011010: dataA <= 32'b10101011011000010010001010000101;
11'b01100011011: dataA <= 32'b00000001111000101010111011000100;
11'b01100011100: dataA <= 32'b01001111001110110011001001110001;
11'b01100011101: dataA <= 32'b00001110101100111101000110110001;
11'b01100011110: dataA <= 32'b00111011010110000110101100110100;
11'b01100011111: dataA <= 32'b00000101000010010000100010111101;
11'b01100100000: dataA <= 32'b00011101100100110001000110001001;
11'b01100100001: dataA <= 32'b00001001111110011101111010001101;
11'b01100100010: dataA <= 32'b01100110101100001011011000101101;
11'b01100100011: dataA <= 32'b00001101101010011111010001110011;
11'b01100100100: dataA <= 32'b10110000101100011001110101001001;
11'b01100100101: dataA <= 32'b00001000111011111101001001110100;
11'b01100100110: dataA <= 32'b00110110011000100100001100000100;
11'b01100100111: dataA <= 32'b00001001001001001111000101100100;
11'b01100101000: dataA <= 32'b01000111011110111011110101011110;
11'b01100101001: dataA <= 32'b00000111100111101000011010101010;
11'b01100101010: dataA <= 32'b10110101011001000010100010101110;
11'b01100101011: dataA <= 32'b00000101011001011001111010110100;
11'b01100101100: dataA <= 32'b10010101110110101001001001001001;
11'b01100101101: dataA <= 32'b00000011001110011110101101110110;
11'b01100101110: dataA <= 32'b11111010110011011100101111010000;
11'b01100101111: dataA <= 32'b00001010100010100100010010100100;
11'b01100110000: dataA <= 32'b01011100001110011011101000010010;
11'b01100110001: dataA <= 32'b00001000010111111011011010000000;
11'b01100110010: dataA <= 32'b10010101001111101011000100111101;
11'b01100110011: dataA <= 32'b00000100110011011101000100010101;
11'b01100110100: dataA <= 32'b10110000111110100100000101111001;
11'b01100110101: dataA <= 32'b00000101101001010000110111101010;
11'b01100110110: dataA <= 32'b11100101000001110001110110001101;
11'b01100110111: dataA <= 32'b00000000101101110110011011001001;
11'b01100111000: dataA <= 32'b01001110110001111100011110001011;
11'b01100111001: dataA <= 32'b00001001100111011110101110000000;
11'b01100111010: dataA <= 32'b01010111110010011101101011110011;
11'b01100111011: dataA <= 32'b00001110110111100101111011010100;
11'b01100111100: dataA <= 32'b10110110011010001001000111000111;
11'b01100111101: dataA <= 32'b00001001111001101111100001000100;
11'b01100111110: dataA <= 32'b01101110110000100110011101101010;
11'b01100111111: dataA <= 32'b00001101111001111101010001000101;
11'b01101000000: dataA <= 32'b00011011011010010100111111010000;
11'b01101000001: dataA <= 32'b00001011001101001101101111001011;
11'b01101000010: dataA <= 32'b10100000011100011001110000101101;
11'b01101000011: dataA <= 32'b00000101010011001001100101001000;
11'b01101000100: dataA <= 32'b11100001100111001100001010110100;
11'b01101000101: dataA <= 32'b00000111010110100111001111010011;
11'b01101000110: dataA <= 32'b10100110011101011001110000110000;
11'b01101000111: dataA <= 32'b00001101000111001111011010001000;
11'b01101001000: dataA <= 32'b10110010011101111001001010000011;
11'b01101001001: dataA <= 32'b00000111100001101100001010011010;
11'b01101001010: dataA <= 32'b00100001010010110000100001010101;
11'b01101001011: dataA <= 32'b00001010100010110000010010100100;
11'b01101001100: dataA <= 32'b00011000111010010101011011111100;
11'b01101001101: dataA <= 32'b00000111011101111011001010100010;
11'b01101001110: dataA <= 32'b10001100111110000000100010101011;
11'b01101001111: dataA <= 32'b00000111110111010111101110111000;
11'b01101010000: dataA <= 32'b01011000110110001110001011010101;
11'b01101010001: dataA <= 32'b00000010110011100110101100001011;
11'b01101010010: dataA <= 32'b00101100011001100101011000110010;
11'b01101010011: dataA <= 32'b00000111001110100100110000001101;
11'b01101010100: dataA <= 32'b01100000111110100000010110001011;
11'b01101010101: dataA <= 32'b00001011010110101001110001100100;
11'b01101010110: dataA <= 32'b00101010110110101010000100110010;
11'b01101010111: dataA <= 32'b00000101100101001100101110001100;
11'b01101011000: dataA <= 32'b11101111101001001011111001101010;
11'b01101011001: dataA <= 32'b00000000101010001101000010001110;
11'b01101011010: dataA <= 32'b10100000010000100001100100101011;
11'b01101011011: dataA <= 32'b00000100100010011000101001100001;
11'b01101011100: dataA <= 32'b01010110111100101011110101101001;
11'b01101011101: dataA <= 32'b00001010110110101001110110010000;
11'b01101011110: dataA <= 32'b11111100110110011011011011101000;
11'b01101011111: dataA <= 32'b00001111010000111001010011101011;
11'b01101100000: dataA <= 32'b01101100111000001011000011010001;
11'b01101100001: dataA <= 32'b00001110110101110011100010010100;
11'b01101100010: dataA <= 32'b10011100000110111010111110001000;
11'b01101100011: dataA <= 32'b00000101101110010001001101000000;
11'b01101100100: dataA <= 32'b00100011111010110010000101111010;
11'b01101100101: dataA <= 32'b00001010110000101001011010001111;
11'b01101100110: dataA <= 32'b01011110111101010010110111101000;
11'b01101100111: dataA <= 32'b00000111000001000101010001111010;
11'b01101101000: dataA <= 32'b10001101011011011010111100110000;
11'b01101101001: dataA <= 32'b00001011000100101000100100010101;
11'b01101101010: dataA <= 32'b01010101011100011100000001010111;
11'b01101101011: dataA <= 32'b00000110000001011000011101101100;
11'b01101101100: dataA <= 32'b00101101110100110001000110000010;
11'b01101101101: dataA <= 32'b00001100010001110101011111101010;
11'b01101101110: dataA <= 32'b10100000101101000100101001100110;
11'b01101101111: dataA <= 32'b00001100011011110101011110011001;
11'b01101110000: dataA <= 32'b10110001010000001011101000000100;
11'b01101110001: dataA <= 32'b00000011111100101000110011001011;
11'b01101110010: dataA <= 32'b00010011011010100010101001110000;
11'b01101110011: dataA <= 32'b00001101100111111100101110001001;
11'b01101110100: dataA <= 32'b01111101000010100110011101010000;
11'b01101110101: dataA <= 32'b00000010100101001100110011000100;
11'b01101110110: dataA <= 32'b11100101100000010010010101001011;
11'b01101110111: dataA <= 32'b00001100111011101001111010011100;
11'b01101111000: dataA <= 32'b10100010100100001100101000001100;
11'b01101111001: dataA <= 32'b00001100000110100011010001101011;
11'b01101111010: dataA <= 32'b11101010100100001011000011101011;
11'b01101111011: dataA <= 32'b00001010111001111100110101111100;
11'b01101111100: dataA <= 32'b01101100001000101101001001100010;
11'b01101111101: dataA <= 32'b00001000001000010011010001100100;
11'b01101111110: dataA <= 32'b00001101101110110011011000011110;
11'b01101111111: dataA <= 32'b00000110001000100000010110010010;
11'b01110000000: dataA <= 32'b00110111000100110011010010110010;
11'b01110000001: dataA <= 32'b00000111011011100101111010111100;
11'b01110000010: dataA <= 32'b10011111111010001000111000001000;
11'b01110000011: dataA <= 32'b00000011110010011010110010010110;
11'b01110000100: dataA <= 32'b01110110011111011011011110101010;
11'b01110000101: dataA <= 32'b00000111100001011010010010101100;
11'b01110000110: dataA <= 32'b01010100010010011011011000110001;
11'b01110000111: dataA <= 32'b00001001010110111101000001010000;
11'b01110001000: dataA <= 32'b11011001010111011001110111111110;
11'b01110001001: dataA <= 32'b00000101110101011111001000110110;
11'b01110001010: dataA <= 32'b01101110110010100011110111111010;
11'b01110001011: dataA <= 32'b00000100101011010001000011010001;
11'b01110001100: dataA <= 32'b00100100111101011010000110001110;
11'b01110001101: dataA <= 32'b00000000110010101100001010101001;
11'b01110001110: dataA <= 32'b01001111000010000100011100100110;
11'b01110001111: dataA <= 32'b00000111100111011010110001010000;
11'b01110010000: dataA <= 32'b01100001110110101101001100010000;
11'b01110010001: dataA <= 32'b00001111010001101111110011010011;
11'b01110010010: dataA <= 32'b01101100001001100001000101101001;
11'b01110010011: dataA <= 32'b00001011011000110101010001001101;
11'b01110010100: dataA <= 32'b11101010100101000111001100000110;
11'b01110010101: dataA <= 32'b00001111010011111100111001010101;
11'b01110010110: dataA <= 32'b01011111011110011100101110101010;
11'b01110010111: dataA <= 32'b00001010101011010111111011000010;
11'b01110011000: dataA <= 32'b10011000011100001011000000110010;
11'b01110011001: dataA <= 32'b00000110010101010001110000100001;
11'b01110011010: dataA <= 32'b11100111100011001011001011010010;
11'b01110011011: dataA <= 32'b00001000010110101001000111001010;
11'b01110011100: dataA <= 32'b10100000011001000010010001010110;
11'b01110011101: dataA <= 32'b00001011000100010101100101100000;
11'b01110011110: dataA <= 32'b01101010010001011001010111100010;
11'b01110011111: dataA <= 32'b00000100100010100010000110000010;
11'b01110100000: dataA <= 32'b11100101001110000000010010111010;
11'b01110100001: dataA <= 32'b00001000000001100110001010100011;
11'b01110100010: dataA <= 32'b11011000111110100101001101111001;
11'b01110100011: dataA <= 32'b00001001111101111010110110001001;
11'b01110100100: dataA <= 32'b01001101001101011000110010001111;
11'b01110100101: dataA <= 32'b00001001010111100001110010001000;
11'b01110100110: dataA <= 32'b10010110111110100101101011110010;
11'b01110100111: dataA <= 32'b00000011110111100010101000001100;
11'b01110101000: dataA <= 32'b01100100010001111101101001010001;
11'b01110101001: dataA <= 32'b00000110101111100000101100100110;
11'b01110101010: dataA <= 32'b10100000111101110000010101101100;
11'b01110101011: dataA <= 32'b00001100010011110011100101100100;
11'b01110101100: dataA <= 32'b11101000101110010001100101010100;
11'b01110101101: dataA <= 32'b00000011101000001010111110001011;
11'b01110101110: dataA <= 32'b01110101011101001100011000001001;
11'b01110101111: dataA <= 32'b00000000110000001111001110101110;
11'b01110110000: dataA <= 32'b00011000010100001010110100001110;
11'b01110110001: dataA <= 32'b00000010000110010100110001000010;
11'b01110110010: dataA <= 32'b01010111000100110100110100001011;
11'b01110110011: dataA <= 32'b00001011110011110011101001100000;
11'b01110110100: dataA <= 32'b10111000011110010011001001100110;
11'b01110110101: dataA <= 32'b00001111001010111010111111100010;
11'b01110110110: dataA <= 32'b00101000101100001100100011110101;
11'b01110110111: dataA <= 32'b00001111001111111001010010010100;
11'b01110111000: dataA <= 32'b10010000001010101010001100000100;
11'b01110111001: dataA <= 32'b00000101010000010101011000100001;
11'b01110111010: dataA <= 32'b11101111110110010001100111111011;
11'b01110111011: dataA <= 32'b00001010101110101101010010101110;
11'b01110111100: dataA <= 32'b10011110111101001011010110001001;
11'b01110111101: dataA <= 32'b00000100000010001011100101101010;
11'b01110111110: dataA <= 32'b11010011101011000001111100001100;
11'b01110111111: dataA <= 32'b00001000100011100010100000101110;
11'b01111000000: dataA <= 32'b10011101100000100101000011011011;
11'b01111000001: dataA <= 32'b00000011100100010100100101110100;
11'b01111000010: dataA <= 32'b00110101101000010010010011100101;
11'b01111000011: dataA <= 32'b00001100001101111001001011001001;
11'b01111000100: dataA <= 32'b01011100101101001101000111100101;
11'b01111000101: dataA <= 32'b00001101110111111001001001111001;
11'b01111000110: dataA <= 32'b11110011000000001101000110000101;
11'b01111000111: dataA <= 32'b00000110111110100100101111000010;
11'b01111001000: dataA <= 32'b00011001100010010010011001101110;
11'b01111001001: dataA <= 32'b00001011100100110110011001101001;
11'b01111001010: dataA <= 32'b01111010101010111101111100101011;
11'b01111001011: dataA <= 32'b00000001001010001011000011000011;
11'b01111001100: dataA <= 32'b01101011011100001011110100101101;
11'b01111001101: dataA <= 32'b00001110110111110011101110100100;
11'b01111001110: dataA <= 32'b11011110100100011110000111101100;
11'b01111001111: dataA <= 32'b00001010000011100111001101101011;
11'b01111010000: dataA <= 32'b11100100011100001100100011001111;
11'b01111010001: dataA <= 32'b00001100010110111000011110000100;
11'b01111010010: dataA <= 32'b10100000000101000110000110100010;
11'b01111010011: dataA <= 32'b00000110101001010111011101101100;
11'b01111010100: dataA <= 32'b11011001111010101010101011011101;
11'b01111010101: dataA <= 32'b00000100101010010110011001111001;
11'b01111010110: dataA <= 32'b01110110110100110100010011110110;
11'b01111010111: dataA <= 32'b00001001011010101111110010110011;
11'b01111011000: dataA <= 32'b00101011110101100001000110101001;
11'b01111011001: dataA <= 32'b00000100010101011000110110110110;
11'b01111011010: dataA <= 32'b11101110010011001010011101000101;
11'b01111011011: dataA <= 32'b00000101000010010010011010101011;
11'b01111011100: dataA <= 32'b00001100011110001011001000110001;
11'b01111011101: dataA <= 32'b00001010110101111100101000101001;
11'b01111011110: dataA <= 32'b10011101011010111001001010111110;
11'b01111011111: dataA <= 32'b00000110110110100001001001011111;
11'b01111100000: dataA <= 32'b10101010100110011011011001111001;
11'b01111100001: dataA <= 32'b00000100001110010011001110101000;
11'b01111100010: dataA <= 32'b10100100111001000010100101110000;
11'b01111100011: dataA <= 32'b00000001111000100000000110000000;
11'b01111100100: dataA <= 32'b00010001001110000100011010100011;
11'b01111100101: dataA <= 32'b00000110001000011000110100101001;
11'b01111100110: dataA <= 32'b01101011110010110100101011101101;
11'b01111100111: dataA <= 32'b00001111001011110111100011000010;
11'b01111101000: dataA <= 32'b11100000000101000001100100001011;
11'b01111101001: dataA <= 32'b00001100110100110111000001100101;
11'b01111101010: dataA <= 32'b00100100100001110111101010000011;
11'b01111101011: dataA <= 32'b00001111001110111010100001110110;
11'b01111101100: dataA <= 32'b10100101011010011100001101000101;
11'b01111101101: dataA <= 32'b00001001101001100001111010100001;
11'b01111101110: dataA <= 32'b11010100100100001100100001111000;
11'b01111101111: dataA <= 32'b00000111010110011101111000001010;
11'b01111110000: dataA <= 32'b00101101011010111010011011101111;
11'b01111110001: dataA <= 32'b00001001010101101010111110111010;
11'b01111110010: dataA <= 32'b01011000011100110011010010111011;
11'b01111110011: dataA <= 32'b00001000100011011101101000111001;
11'b01111110100: dataA <= 32'b01100000001000111010000101000011;
11'b01111110101: dataA <= 32'b00000010000101010110000101110010;
11'b01111110110: dataA <= 32'b01100111001001010000010101011101;
11'b01111110111: dataA <= 32'b00000101000010011010001010011011;
11'b01111111000: dataA <= 32'b11011001000110101100101111010011;
11'b01111111001: dataA <= 32'b00001100011010110110100001101001;
11'b01111111010: dataA <= 32'b01010001011000110001100010110011;
11'b01111111011: dataA <= 32'b00001010010110101001101101011000;
11'b01111111100: dataA <= 32'b00010111000110111101001100001111;
11'b01111111101: dataA <= 32'b00000101011010011110101000011110;
11'b01111111110: dataA <= 32'b01011100010010001101101001010000;
11'b01111111111: dataA <= 32'b00000110110000011100101101001111;
11'b10000000000: dataA <= 32'b11100000111101000000100101001110;
11'b10000000001: dataA <= 32'b00001100101111111001010101110100;
11'b10000000010: dataA <= 32'b11100100101001110001100110010110;
11'b10000000011: dataA <= 32'b00000010101011001101001110001011;
11'b10000000100: dataA <= 32'b10111001001001011101000111001001;
11'b10000000101: dataA <= 32'b00000001010110010011011011000101;
11'b10000000110: dataA <= 32'b00010000011100001100000100010001;
11'b10000000111: dataA <= 32'b00000000101011010010111000110011;
11'b10000001000: dataA <= 32'b11100011010010011110010101110111;
11'b10000001001: dataA <= 32'b00001001101000110100011000001100;
11'b10000001010: dataA <= 32'b11001110001101100011010011001100;
11'b10000001011: dataA <= 32'b00000101000001011110001001010000;
11'b10000001100: dataA <= 32'b01010110101110010111101010111000;
11'b10000001101: dataA <= 32'b00000111100001101000001110000011;
11'b10000001110: dataA <= 32'b11000101011101000010100010000111;
11'b10000001111: dataA <= 32'b00001000010101101101010100110110;
11'b10000010000: dataA <= 32'b10111010100000110011011101110000;
11'b10000010001: dataA <= 32'b00000111001010101000100111011010;
11'b10000010010: dataA <= 32'b10011111000001101101100100110011;
11'b10000010011: dataA <= 32'b00000001010111110011101001010100;
11'b10000010100: dataA <= 32'b10110101011000111001110110000111;
11'b10000010101: dataA <= 32'b00000001101110010000111011011110;
11'b10000010110: dataA <= 32'b01110001000110100110111101111001;
11'b10000010111: dataA <= 32'b00000010011000010011010110010100;
11'b10000011000: dataA <= 32'b10110100010101001111010010111000;
11'b10000011001: dataA <= 32'b00000110100111100100001100100001;
11'b10000011010: dataA <= 32'b00010111000110100101100010110000;
11'b10000011011: dataA <= 32'b00001011100100100100001100101100;
11'b10000011100: dataA <= 32'b11100000011010100111100010110011;
11'b10000011101: dataA <= 32'b00001111010010010110110101011001;
11'b10000011110: dataA <= 32'b10110001001101001011010111001100;
11'b10000011111: dataA <= 32'b00000010001000001100010000100100;
11'b10000100000: dataA <= 32'b11010100001010111010000101100110;
11'b10000100001: dataA <= 32'b00000101011101100001101001101001;
11'b10000100010: dataA <= 32'b11101110101001111111100110110110;
11'b10000100011: dataA <= 32'b00001011100010110110011010001010;
11'b10000100100: dataA <= 32'b10010011000011000111000110010000;
11'b10000100101: dataA <= 32'b00000001101011100110110001111100;
11'b10000100110: dataA <= 32'b11001110110110010111100111111001;
11'b10000100111: dataA <= 32'b00001011000111001110001110011011;
11'b10000101000: dataA <= 32'b10000010111111000101110001010010;
11'b10000101001: dataA <= 32'b00000100110010101111010010010100;
11'b10000101010: dataA <= 32'b00111101001101010010101110101001;
11'b10000101011: dataA <= 32'b00000101010110001101010000111100;
11'b10000101100: dataA <= 32'b01011010010010001110011011011000;
11'b10000101101: dataA <= 32'b00001101001101111000100001101010;
11'b10000101110: dataA <= 32'b01111010101000100100110100110010;
11'b10000101111: dataA <= 32'b00001010110111011011001111000010;
11'b10000110000: dataA <= 32'b10001000100001001001100010100101;
11'b10000110001: dataA <= 32'b00000001010101001101011001111010;
11'b10000110010: dataA <= 32'b10001111100101100011101000101110;
11'b10000110011: dataA <= 32'b00001010101010010100000100100110;
11'b10000110100: dataA <= 32'b00101101000100100010001111001010;
11'b10000110101: dataA <= 32'b00001011010010100100111111110101;
11'b10000110110: dataA <= 32'b10010010101001101011001100101100;
11'b10000110111: dataA <= 32'b00000111010111100111011000010010;
11'b10000111000: dataA <= 32'b11011100110101010101111000010100;
11'b10000111001: dataA <= 32'b00001100011100000010111100010011;
11'b10000111010: dataA <= 32'b10100111011110001011110001101010;
11'b10000111011: dataA <= 32'b00000100010011011011001100100110;
11'b10000111100: dataA <= 32'b11111000101010010010010110101000;
11'b10000111101: dataA <= 32'b00000101100001110000010001001001;
11'b10000111110: dataA <= 32'b11000010111100110101110101110111;
11'b10000111111: dataA <= 32'b00001010000110100000010010111100;
11'b10001000000: dataA <= 32'b01010000110111110100010001101011;
11'b10001000001: dataA <= 32'b00000111000001010000001011000100;
11'b10001000010: dataA <= 32'b11101100110110000011000010100101;
11'b10001000011: dataA <= 32'b00000100101100111100111100110010;
11'b10001000100: dataA <= 32'b10010011010110010111101100011100;
11'b10001000101: dataA <= 32'b00001011010001111101000101011111;
11'b10001000110: dataA <= 32'b00101100100101001010000111101000;
11'b10001000111: dataA <= 32'b00001010101101011110101001000010;
11'b10001001000: dataA <= 32'b00001111001101101110011101111010;
11'b10001001001: dataA <= 32'b00000001101110110101000100101110;
11'b10001001010: dataA <= 32'b01000100111101000110000001110101;
11'b10001001011: dataA <= 32'b00000010111011000011010001001100;
11'b10001001100: dataA <= 32'b00100100110000001101011110110101;
11'b10001001101: dataA <= 32'b00000001010101000101001001101011;
11'b10001001110: dataA <= 32'b10100011001110010010101001100001;
11'b10001001111: dataA <= 32'b00001101000111010000010000111100;
11'b10001010000: dataA <= 32'b00101101011100110110011001111010;
11'b10001010001: dataA <= 32'b00001011001011110110101100001101;
11'b10001010010: dataA <= 32'b00100011010010100010000111100111;
11'b10001010011: dataA <= 32'b00001101010101010101000011000111;
11'b10001010100: dataA <= 32'b10001001000110110011101000001101;
11'b10001010101: dataA <= 32'b00001000010010010111000111101101;
11'b10001010110: dataA <= 32'b01011110111100010101110111010101;
11'b10001010111: dataA <= 32'b00000111100110101010001110011100;
11'b10001011000: dataA <= 32'b10010100110100110100011011010011;
11'b10001011001: dataA <= 32'b00000101111010100111100101111011;
11'b10001011010: dataA <= 32'b11100100001110100101000100110001;
11'b10001011011: dataA <= 32'b00001011011101101101011010110001;
11'b10001011100: dataA <= 32'b01001111011110000111101000110111;
11'b10001011101: dataA <= 32'b00000101111110011101011001100110;
11'b10001011110: dataA <= 32'b01011111010001111110100100110100;
11'b10001011111: dataA <= 32'b00001011001010111010101100001011;
11'b10001100000: dataA <= 32'b10011010000101101011000100001000;
11'b10001100001: dataA <= 32'b00001000000001101000001101111000;
11'b10001100010: dataA <= 32'b01011100100101100111101000111001;
11'b10001100011: dataA <= 32'b00001010100010110000011010001011;
11'b10001100100: dataA <= 32'b11000011000101011010000100000011;
11'b10001100101: dataA <= 32'b00000111010100100111011100010101;
11'b10001100110: dataA <= 32'b10111100111001000010011101010100;
11'b10001100111: dataA <= 32'b00001000001010101100101111100011;
11'b10001101000: dataA <= 32'b00011111000001011101010100010000;
11'b10001101001: dataA <= 32'b00000000110001101001110101001100;
11'b10001101010: dataA <= 32'b01101101100101011001001000000110;
11'b10001101011: dataA <= 32'b00000010001001010010101110110111;
11'b10001101100: dataA <= 32'b10101111010110000111001011111101;
11'b10001101101: dataA <= 32'b00000000110011001111001110001100;
11'b10001101110: dataA <= 32'b10111010100100100110010001010011;
11'b10001101111: dataA <= 32'b00001000100111101110010101000000;
11'b10001110000: dataA <= 32'b00010110111110010101110011001100;
11'b10001110001: dataA <= 32'b00001101100111101110010100110011;
11'b10001110010: dataA <= 32'b10101000011101110111100010001111;
11'b10001110011: dataA <= 32'b00001110011000011000101101110001;
11'b10001110100: dataA <= 32'b10101101011001010010111000001100;
11'b10001110101: dataA <= 32'b00000011100100010110000100100011;
11'b10001110110: dataA <= 32'b11100000000111001010111000000101;
11'b10001110111: dataA <= 32'b00000010111010011001100110001001;
11'b10001111000: dataA <= 32'b00110000110101001111010101110101;
11'b10001111001: dataA <= 32'b00001101100110111100101110011011;
11'b10001111010: dataA <= 32'b10010010111010010111100110001111;
11'b10001111011: dataA <= 32'b00000011000111101000111001110100;
11'b10001111100: dataA <= 32'b00010010101001100111100101111000;
11'b10001111101: dataA <= 32'b00001100101010011010000110011100;
11'b10001111110: dataA <= 32'b11000100100110100110100001001100;
11'b10001111111: dataA <= 32'b00000100001111101001011010001100;
11'b10010000000: dataA <= 32'b01110111100101101010011111001111;
11'b10010000001: dataA <= 32'b00000100010011001010111101000011;
11'b10010000010: dataA <= 32'b00100010010001101110011001011010;
11'b10010000011: dataA <= 32'b00001101110001111100110110000010;
11'b10010000100: dataA <= 32'b01111101000000011011100100001111;
11'b10010000101: dataA <= 32'b00001001011000011001001011010011;
11'b10010000110: dataA <= 32'b10001110010001101001000101000010;
11'b10010000111: dataA <= 32'b00000000110000001001001010001010;
11'b10010001000: dataA <= 32'b01001001010101101011001000101110;
11'b10010001001: dataA <= 32'b00001011001101100000000100001101;
11'b10010001010: dataA <= 32'b01101011001100111001001111010000;
11'b10010001011: dataA <= 32'b00001010110100100101000011011110;
11'b10010001100: dataA <= 32'b01011000100001111010111101010000;
11'b10010001101: dataA <= 32'b00000101110110100001011100101001;
11'b10010001110: dataA <= 32'b10011110110101000101000111010011;
11'b10010001111: dataA <= 32'b00001001011110000100100100100010;
11'b10010010000: dataA <= 32'b01100001100010001011110011000110;
11'b10010010001: dataA <= 32'b00000011110000011001001000001101;
11'b10010010010: dataA <= 32'b01111010111110100010101000000111;
11'b10010010011: dataA <= 32'b00001000100001111000100001101001;
11'b10010010100: dataA <= 32'b10000100100100100100110100110100;
11'b10010010101: dataA <= 32'b00001100001001101000010110101101;
11'b10010010110: dataA <= 32'b01010010101011100101110011000111;
11'b10010010111: dataA <= 32'b00001001100001011100000110111101;
11'b10010011000: dataA <= 32'b11101111000010010011000101000010;
11'b10010011001: dataA <= 32'b00000101101010111101010001001001;
11'b10010011010: dataA <= 32'b11001111001101100111101001011110;
11'b10010011011: dataA <= 32'b00001010110011111001011100110110;
11'b10010011100: dataA <= 32'b10110000110001100001101001001001;
11'b10010011101: dataA <= 32'b00001011001111100010101101011001;
11'b10010011110: dataA <= 32'b11001100111101001101111011011101;
11'b10010011111: dataA <= 32'b00000010001001110011010100010100;
11'b10010100000: dataA <= 32'b11001000101000101101000001010000;
11'b10010100001: dataA <= 32'b00000001010110000010111001001011;
11'b10010100010: dataA <= 32'b11100110110100001011111101011010;
11'b10010100011: dataA <= 32'b00000000101111000100110001111010;
11'b10010100100: dataA <= 32'b10011111001110100010111100100100;
11'b10010100101: dataA <= 32'b00001110101100011010001000111011;
11'b10010100110: dataA <= 32'b10100111100100011101000111111011;
11'b10010100111: dataA <= 32'b00001011101101111000111100001011;
11'b10010101000: dataA <= 32'b10011111010010110010111001001000;
11'b10010101001: dataA <= 32'b00001011111000010100111010010111;
11'b10010101010: dataA <= 32'b11001000110110110100001000101101;
11'b10010101011: dataA <= 32'b00000111110010010110111111001110;
11'b10010101100: dataA <= 32'b11011110111100001100010110010100;
11'b10010101101: dataA <= 32'b00001001100111110010011010010100;
11'b10010101110: dataA <= 32'b10010110101100110011011010010101;
11'b10010101111: dataA <= 32'b00000100011000011111101001111011;
11'b10010110000: dataA <= 32'b10101110010110001101100100101111;
11'b10010110001: dataA <= 32'b00001000011110100111100011001010;
11'b10010110010: dataA <= 32'b11001011001101011111100111010111;
11'b10010110011: dataA <= 32'b00000011011011011001010101000101;
11'b10010110100: dataA <= 32'b00011011001101011110010011110001;
11'b10010110101: dataA <= 32'b00001011101101111101000100011010;
11'b10010110110: dataA <= 32'b11100100000101111010110110000110;
11'b10010110111: dataA <= 32'b00001011000010110010011010100000;
11'b10010111000: dataA <= 32'b10100000100100111111000111011001;
11'b10010111001: dataA <= 32'b00001101000101110110101010010011;
11'b10010111010: dataA <= 32'b01000010101101110001110110100001;
11'b10010111011: dataA <= 32'b00000110010011100001100000001100;
11'b10010111100: dataA <= 32'b11111101001101011001111011111000;
11'b10010111101: dataA <= 32'b00001001001010101110111011100100;
11'b10010111110: dataA <= 32'b10011111000001001100110100001101;
11'b10010111111: dataA <= 32'b00000000101011011101111001001011;
11'b10011000000: dataA <= 32'b10100101101110000000111001100111;
11'b10011000001: dataA <= 32'b00000011100101010110100110000111;
11'b10011000010: dataA <= 32'b11101011011101011110111000111110;
11'b10011000011: dataA <= 32'b00000000101101001110111110000100;
11'b10011000100: dataA <= 32'b01111100111100001101000001001110;
11'b10011000101: dataA <= 32'b00001010001000110100100001110000;
11'b10011000110: dataA <= 32'b01011000110101111101110011101001;
11'b10011000111: dataA <= 32'b00001110101100110100100000111010;
11'b10011001000: dataA <= 32'b11101100101001000111010010101011;
11'b10011001001: dataA <= 32'b00001100011100011100101010010001;
11'b10011001010: dataA <= 32'b01100111100001100010011000101100;
11'b10011001011: dataA <= 32'b00000110000010100010000100101010;
11'b10011001100: dataA <= 32'b00101010001011010011111010000110;
11'b10011001101: dataA <= 32'b00000001010101010001011110100010;
11'b10011001110: dataA <= 32'b10110011000100100110010100110011;
11'b10011001111: dataA <= 32'b00001111001100111101000110100011;
11'b10011010000: dataA <= 32'b01010110110001101111100110101110;
11'b10011010001: dataA <= 32'b00000101000100101001000001101100;
11'b10011010010: dataA <= 32'b01010110011100111111000100110101;
11'b10011010011: dataA <= 32'b00001101101110100100000110010100;
11'b10011010100: dataA <= 32'b11001100010010000110110010000111;
11'b10011010101: dataA <= 32'b00000100101101100011100010000100;
11'b10011010110: dataA <= 32'b10101111110001111010001111010101;
11'b10011010111: dataA <= 32'b00000011110000001100101101001010;
11'b10011011000: dataA <= 32'b01101100010101010101110111011010;
11'b10011011001: dataA <= 32'b00001100110101111101001110010010;
11'b10011011010: dataA <= 32'b01111011010100100010100100101101;
11'b10011011011: dataA <= 32'b00000111011001010111000011010100;
11'b10011011100: dataA <= 32'b11011000001010010001001000000001;
11'b10011011101: dataA <= 32'b00000001001010001000110110011010;
11'b10011011110: dataA <= 32'b11000111000101110011001001001111;
11'b10011011111: dataA <= 32'b00001011101111101100001000001011;
11'b10011100000: dataA <= 32'b01100111010101100000101110110110;
11'b10011100001: dataA <= 32'b00001001110110100011000110110111;
11'b10011100010: dataA <= 32'b10011110011110000010111100110100;
11'b10011100011: dataA <= 32'b00000100110100011011011101010000;
11'b10011100100: dataA <= 32'b10100000110100111100010110110011;
11'b10011100101: dataA <= 32'b00000110111110001100010000111001;
11'b10011100110: dataA <= 32'b11011001100010001100000101100011;
11'b10011100111: dataA <= 32'b00000011101100010111000000001011;
11'b10011101000: dataA <= 32'b01111001010010110011001001101000;
11'b10011101001: dataA <= 32'b00001011100010111100110110001001;
11'b10011101010: dataA <= 32'b11001100010000100011100011110001;
11'b10011101011: dataA <= 32'b00001100101100110000100010010101;
11'b10011101100: dataA <= 32'b11011000100011001110110101000100;
11'b10011101101: dataA <= 32'b00001100100100101000000110101101;
11'b10011101110: dataA <= 32'b10101101001010011011011000000001;
11'b10011101111: dataA <= 32'b00000110101001110111100101100001;
11'b10011110000: dataA <= 32'b10001110111100111111000110111110;
11'b10011110001: dataA <= 32'b00001001110101110011101100010101;
11'b10011110010: dataA <= 32'b01110010111110000001101010001010;
11'b10011110011: dataA <= 32'b00001011010001100110110001111001;
11'b10011110100: dataA <= 32'b10001110110000111101001000011110;
11'b10011110101: dataA <= 32'b00000011100101101101100000010011;
11'b10011110110: dataA <= 32'b00001110011000100100000001101011;
11'b10011110111: dataA <= 32'b00000000110000000100100101010011;
11'b10011111000: dataA <= 32'b11101000111100010010011010111101;
11'b10011111001: dataA <= 32'b00000001001010001000011110000010;
11'b10011111010: dataA <= 32'b11011101001110101011011110001000;
11'b10011111011: dataA <= 32'b00001110110001100100001001000010;
11'b10011111100: dataA <= 32'b00011111100100010011110101111010;
11'b10011111101: dataA <= 32'b00001011110000110111010000010010;
11'b10011111110: dataA <= 32'b10011011001111000011101010101001;
11'b10011111111: dataA <= 32'b00001001111010010110110001101111;
11'b10100000000: dataA <= 32'b10001100100110101100111001001110;
11'b10100000001: dataA <= 32'b00000111010001011000110110100111;
11'b10100000010: dataA <= 32'b11011110111100001010110101110011;
11'b10100000011: dataA <= 32'b00001011001001111000101110001100;
11'b10100000100: dataA <= 32'b10011010101001000010101001010110;
11'b10100000101: dataA <= 32'b00000010110100010111100110000011;
11'b10100000110: dataA <= 32'b10110100100001111101100101001100;
11'b10100000111: dataA <= 32'b00000101011110100001100111011011;
11'b10100001000: dataA <= 32'b11001000111100110110110101110110;
11'b10100001001: dataA <= 32'b00000001010110010101001100110100;
11'b10100001010: dataA <= 32'b11011001001001000101100011101110;
11'b10100001011: dataA <= 32'b00001100010000111001011000111000;
11'b10100001100: dataA <= 32'b10110000001110001010111000000101;
11'b10100001101: dataA <= 32'b00001101100101111000101011001001;
11'b10100001110: dataA <= 32'b11100100101000011110000101011000;
11'b10100001111: dataA <= 32'b00001110101010111010111110010011;
11'b10100010000: dataA <= 32'b11001000011010010001111001100010;
11'b10100010001: dataA <= 32'b00000101110001011011011100001010;
11'b10100010010: dataA <= 32'b00110111100101111001011010011010;
11'b10100010011: dataA <= 32'b00001010001100101111000111001110;
11'b10100010100: dataA <= 32'b11011111000001000100000100101011;
11'b10100010101: dataA <= 32'b00000010000110010011110001011010;
11'b10100010110: dataA <= 32'b10011101101110100001001011001001;
11'b10100010111: dataA <= 32'b00000110000011011100100001010111;
11'b10100011000: dataA <= 32'b11100011100000111110000101111110;
11'b10100011001: dataA <= 32'b00000001101000010000110001111100;
11'b10100011010: dataA <= 32'b01111101010100001011110010001001;
11'b10100011011: dataA <= 32'b00001011101010111000110110100000;
11'b10100011100: dataA <= 32'b10011010110001100101100101100110;
11'b10100011101: dataA <= 32'b00001110110010111000110101011001;
11'b10100011110: dataA <= 32'b00110000110100100110010100000111;
11'b10100011111: dataA <= 32'b00001001011110100000101010101010;
11'b10100100000: dataA <= 32'b10011111100101111010001001001101;
11'b10100100001: dataA <= 32'b00001001000010101110001001000001;
11'b10100100010: dataA <= 32'b10110100010111001101001011101000;
11'b10100100011: dataA <= 32'b00000000101111001101001110111010;
11'b10100100100: dataA <= 32'b00110001010000001101000100010000;
11'b10100100101: dataA <= 32'b00001111010001111011011110101100;
11'b10100100110: dataA <= 32'b00011000101000111111000111001101;
11'b10100100111: dataA <= 32'b00000111100010101001001001101100;
11'b10100101000: dataA <= 32'b10011110011000011110000011110010;
11'b10100101001: dataA <= 32'b00001101010010110000001110001100;
11'b10100101010: dataA <= 32'b11010110000101100110100100000100;
11'b10100101011: dataA <= 32'b00000101001010011101100001110100;
11'b10100101100: dataA <= 32'b00100011111010010010011101111010;
11'b10100101101: dataA <= 32'b00000100001101010000100001100010;
11'b10100101110: dataA <= 32'b10110010100000111101000101011001;
11'b10100101111: dataA <= 32'b00001011011000110111100010101010;
11'b10100110000: dataA <= 32'b01110101101000111001100101001010;
11'b10100110001: dataA <= 32'b00000101111000010110111011001101;
11'b10100110010: dataA <= 32'b01100100001010110001101010100010;
11'b10100110011: dataA <= 32'b00000010100101001100100110100011;
11'b10100110100: dataA <= 32'b01001000110010000010111001010000;
11'b10100110101: dataA <= 32'b00001011010010110110010100010010;
11'b10100110110: dataA <= 32'b10100011011010010000101101011011;
11'b10100110111: dataA <= 32'b00001000010111100011000110000111;
11'b10100111000: dataA <= 32'b01100100100010010011001011010111;
11'b10100111001: dataA <= 32'b00000100010001010111011010000000;
11'b10100111010: dataA <= 32'b11100010110100111011010110010001;
11'b10100111011: dataA <= 32'b00000011111100010110000101011000;
11'b10100111100: dataA <= 32'b01010101011010001100001000000010;
11'b10100111101: dataA <= 32'b00000100101010010110111000010010;
11'b10100111110: dataA <= 32'b10110011100110111011111011001010;
11'b10100111111: dataA <= 32'b00001101100110111011001110101001;
11'b10101000000: dataA <= 32'b00010110000100101010010011101110;
11'b10101000001: dataA <= 32'b00001101010000110100101101111110;
11'b10101000010: dataA <= 32'b00011110011110011111100111100010;
11'b10101000011: dataA <= 32'b00001110101000110010010010001110;
11'b10101000100: dataA <= 32'b01101011010110011011111010100010;
11'b10101000101: dataA <= 32'b00001000001000101101110110000001;
11'b10101000110: dataA <= 32'b00010000110000011110000011111100;
11'b10101000111: dataA <= 32'b00001000110110100111111000001100;
11'b10101001000: dataA <= 32'b10110001001110100001101011001100;
11'b10101001001: dataA <= 32'b00001010010100101000111010100001;
11'b10101001010: dataA <= 32'b01010010100100101100000101011110;
11'b10101001011: dataA <= 32'b00000110000011100111101000100010;
11'b10101001100: dataA <= 32'b10010110001100101011000011000110;
11'b10101001101: dataA <= 32'b00000000101010001100010001011010;
11'b10101001110: dataA <= 32'b00101001000100101001010111111110;
11'b10101001111: dataA <= 32'b00000010100101010000010010010011;
11'b10101010000: dataA <= 32'b00011011001010110011111111001110;
11'b10101010001: dataA <= 32'b00001101110110101110010001010010;
11'b10101010010: dataA <= 32'b00010111100100011010100011110111;
11'b10101010011: dataA <= 32'b00001011010011110001100000110001;
11'b10101010100: dataA <= 32'b00011001001011000100011011101100;
11'b10101010101: dataA <= 32'b00000111111011011010101100111111;
11'b10101010110: dataA <= 32'b10010010010110100101011001001111;
11'b10101010111: dataA <= 32'b00000111010001011010110001111111;
11'b10101011000: dataA <= 32'b00011110111100100001100101010001;
11'b10101011001: dataA <= 32'b00001100001100111011000001111101;
11'b10101011010: dataA <= 32'b10011110100101011001110111110111;
11'b10101011011: dataA <= 32'b00000010010000010001011010000011;
11'b10101011100: dataA <= 32'b10111000110101101101010101101010;
11'b10101011101: dataA <= 32'b00000010111011011001100011010100;
11'b10101011110: dataA <= 32'b11001010101000010101100100110100;
11'b10101011111: dataA <= 32'b00000000110000010011000100101011;
endcase
if (enB)
case(addrB)
11'b00000000000: dataB <= 32'b00100101001110110101110111011000;
11'b00000000001: dataB <= 32'b00001000000111101100001100011110;
11'b00000000010: dataB <= 32'b10000110011101011011100010101111;
11'b00000000011: dataB <= 32'b00000010100100010100001100110001;
11'b00000000100: dataB <= 32'b01010100110111000111001100010101;
11'b00000000101: dataB <= 32'b00000101000010011110001001111011;
11'b00000000110: dataB <= 32'b10001101101100111011010001001100;
11'b00000000111: dataB <= 32'b00001000110100101111001001011111;
11'b00000001000: dataB <= 32'b10110010010000101100001101001011;
11'b00000001001: dataB <= 32'b00000110001011100010100011000001;
11'b00000001010: dataB <= 32'b00100001000010000101110101110110;
11'b00000001011: dataB <= 32'b00000011011011111001011001011101;
11'b00000001100: dataB <= 32'b01110111000100100010110100101001;
11'b00000001101: dataB <= 32'b00000001110011010001000111110101;
11'b00000001110: dataB <= 32'b00110000111011000110001111010100;
11'b00000001111: dataB <= 32'b00000100011100011001011110011100;
11'b00000010000: dataB <= 32'b11101010000101111111100100111011;
11'b00000010001: dataB <= 32'b00000101001000011010001100001010;
11'b00000010010: dataB <= 32'b00011001001010110100110011010100;
11'b00000010011: dataB <= 32'b00001001000010011010001100110101;
11'b00000010100: dataB <= 32'b10011010011111001110110011110111;
11'b00000010101: dataB <= 32'b00001111001101010100111101000010;
11'b00000010110: dataB <= 32'b11110011000001000100000110101101;
11'b00000010111: dataB <= 32'b00000001001101000100100000110101;
11'b00000011000: dataB <= 32'b00001010010110100001100100001000;
11'b00000011001: dataB <= 32'b00000111111110100111100101010010;
11'b00000011010: dataB <= 32'b10101000011110100111101000010111;
11'b00000011011: dataB <= 32'b00001000100001101110001010000010;
11'b00000011100: dataB <= 32'b10010101001111100110000110110001;
11'b00000011101: dataB <= 32'b00000001010000100100101110000100;
11'b00000011110: dataB <= 32'b10001101000011000111001001011000;
11'b00000011111: dataB <= 32'b00001001000101000110011110010011;
11'b00000100000: dataB <= 32'b01000011010011010100110010010111;
11'b00000100001: dataB <= 32'b00000101010101110001000110011100;
11'b00000100010: dataB <= 32'b11111100111001001011011101000100;
11'b00000100011: dataB <= 32'b00000110110111010001011101000100;
11'b00000100100: dataB <= 32'b10010000011010100110001100110101;
11'b00000100101: dataB <= 32'b00001100001001110000010001010010;
11'b00000100110: dataB <= 32'b10110100010100110110000101010101;
11'b00000100111: dataB <= 32'b00001100010100011101010010101001;
11'b00000101000: dataB <= 32'b11000100110100110010010001001010;
11'b00000101001: dataB <= 32'b00000010111010010011100101101010;
11'b00000101010: dataB <= 32'b01011001101101011011111000001101;
11'b00000101011: dataB <= 32'b00001001001001001010010001001111;
11'b00000101100: dataB <= 32'b11101100111000010011011101100101;
11'b00000101101: dataB <= 32'b00001011101111100010111011110011;
11'b00000101110: dataB <= 32'b11010000110101100011011011101001;
11'b00000101111: dataB <= 32'b00001000110111101101010000001011;
11'b00000110000: dataB <= 32'b00011010111001101110001000110011;
11'b00000110001: dataB <= 32'b00001110011000000011010000011101;
11'b00000110010: dataB <= 32'b01101101010110000011100001001111;
11'b00000110011: dataB <= 32'b00000101010110011101010001001111;
11'b00000110100: dataB <= 32'b10110010011001111010000101001001;
11'b00000110101: dataB <= 32'b00000011000100100110001000110010;
11'b00000110110: dataB <= 32'b00000011010001001110100111011000;
11'b00000110111: dataB <= 32'b00001000000101010110010111000100;
11'b00000111000: dataB <= 32'b10001111000011110011000001010000;
11'b00000111001: dataB <= 32'b00000100000010001000011011000011;
11'b00000111010: dataB <= 32'b11101010101001111011000001001010;
11'b00000111011: dataB <= 32'b00000100001111111010100100101011;
11'b00000111100: dataB <= 32'b10011001011111000111001110011000;
11'b00000111101: dataB <= 32'b00001011001110111100110010000111;
11'b00000111110: dataB <= 32'b11100110011100110010110110001001;
11'b00000111111: dataB <= 32'b00001010001011011100101100110010;
11'b00001000000: dataB <= 32'b11010011011010000110101111010101;
11'b00001000001: dataB <= 32'b00000001110011110100110001001110;
11'b00001000010: dataB <= 32'b00000111010001100110100011011001;
11'b00001000011: dataB <= 32'b00000101011110001001100101010101;
11'b00001000100: dataB <= 32'b01100010101100101110101111010000;
11'b00001000101: dataB <= 32'b00000010111010001001011101100011;
11'b00001000110: dataB <= 32'b01100101001001111010010111000001;
11'b00001000111: dataB <= 32'b00001011000100001000100001000101;
11'b00001001000: dataB <= 32'b01110011010001010111001011111000;
11'b00001001001: dataB <= 32'b00001001101001110000011100100110;
11'b00001001010: dataB <= 32'b00100101001110001001110110001000;
11'b00001001011: dataB <= 32'b00001101110000010111001011100110;
11'b00001001100: dataB <= 32'b00001011011010101010110111101101;
11'b00001001101: dataB <= 32'b00001000110001011001001011110100;
11'b00001001110: dataB <= 32'b00011111000000110110111000110101;
11'b00001001111: dataB <= 32'b00000110000111100000001010100100;
11'b00001010000: dataB <= 32'b11010011000000111101001011110000;
11'b00001010001: dataB <= 32'b00001000011011101101011101110011;
11'b00001010010: dataB <= 32'b01011010001110101100100101010100;
11'b00001010011: dataB <= 32'b00001101111010110001001110010001;
11'b00001010100: dataB <= 32'b10010101101010110111011010010110;
11'b00001010101: dataB <= 32'b00001000011110100011011001111110;
11'b00001010110: dataB <= 32'b00100111001011001101001000111000;
11'b00001010111: dataB <= 32'b00000110101000100010000101000111;
11'b00001011000: dataB <= 32'b11000010110101011100000011010011;
11'b00001011001: dataB <= 32'b00000001001001001100011000011010;
11'b00001011010: dataB <= 32'b01010010111111100110001100110001;
11'b00001011011: dataB <= 32'b00000010100101010100010001110011;
11'b00001011100: dataB <= 32'b10010111111000111100010000110010;
11'b00001011101: dataB <= 32'b00001001110011110000111110001111;
11'b00001011110: dataB <= 32'b11100110000100111101001100001000;
11'b00001011111: dataB <= 32'b00000101001101011100100010011000;
11'b00001100000: dataB <= 32'b10100001000010011101100110110111;
11'b00001100001: dataB <= 32'b00000101111110111101000101110101;
11'b00001100010: dataB <= 32'b11110110110100011011110011101100;
11'b00001100011: dataB <= 32'b00000010111000010011010011110011;
11'b00001100100: dataB <= 32'b11101110101011011101001111001110;
11'b00001100101: dataB <= 32'b00000110111110011111100010011011;
11'b00001100110: dataB <= 32'b01011110000110100111100111011101;
11'b00001100111: dataB <= 32'b00000100001011010000010100001100;
11'b00001101000: dataB <= 32'b00011011001110111100000100111000;
11'b00001101001: dataB <= 32'b00000110000010010000010101001110;
11'b00001101010: dataB <= 32'b01010100100111101101110101111010;
11'b00001101011: dataB <= 32'b00001110000111010101000100111011;
11'b00001101100: dataB <= 32'b10110000110001001100110110001110;
11'b00001101101: dataB <= 32'b00000001010011000010111001001110;
11'b00001101110: dataB <= 32'b11000100101001111001010011001011;
11'b00001101111: dataB <= 32'b00001010111101101111011101000010;
11'b00001110000: dataB <= 32'b11100010011011001110111001110110;
11'b00001110001: dataB <= 32'b00000110000001100010000101110010;
11'b00001110010: dataB <= 32'b10011001010011110100100111010010;
11'b00001110011: dataB <= 32'b00000010010101100000101110001100;
11'b00001110100: dataB <= 32'b01001111010011100110001010110110;
11'b00001110101: dataB <= 32'b00000111000100000010110110001011;
11'b00001110110: dataB <= 32'b11001001100111011011110011111011;
11'b00001110111: dataB <= 32'b00000110110110110000111010011011;
11'b00001111000: dataB <= 32'b10111000100001000100001010100001;
11'b00001111001: dataB <= 32'b00001000011000010111100101010101;
11'b00001111010: dataB <= 32'b01001010100110111101011101010001;
11'b00001111011: dataB <= 32'b00001010100110100110000101001011;
11'b00001111100: dataB <= 32'b01101010001001010110110110110110;
11'b00001111101: dataB <= 32'b00001100110001100001010010001001;
11'b00001111110: dataB <= 32'b00000101001100100011010000101111;
11'b00001111111: dataB <= 32'b00000101011101011011101101011011;
11'b00010000000: dataB <= 32'b10100011110001100100010111101101;
11'b00010000001: dataB <= 32'b00000111101000000100100101111111;
11'b00010000010: dataB <= 32'b01101010110000010100111011000010;
11'b00010000011: dataB <= 32'b00001011001100100010111011101010;
11'b00010000100: dataB <= 32'b01001111000001011011111010000110;
11'b00010000101: dataB <= 32'b00001010010110101111001000010101;
11'b00010000110: dataB <= 32'b00011010111110001110001001110010;
11'b00010000111: dataB <= 32'b00001111010010001001100100110110;
11'b00010001000: dataB <= 32'b10110001001110000011100001110100;
11'b00010001001: dataB <= 32'b00000110011000100001010001111111;
11'b00010001010: dataB <= 32'b10101000001101100010010100001100;
11'b00010001011: dataB <= 32'b00000001001000011010000100101011;
11'b00010001100: dataB <= 32'b01001001100101110110111000111000;
11'b00010001101: dataB <= 32'b00000110000110010000011110111011;
11'b00010001110: dataB <= 32'b10010001001111011001100010010101;
11'b00010001111: dataB <= 32'b00000010000110000010101110111010;
11'b00010010000: dataB <= 32'b11100100100101101011000000101111;
11'b00010010001: dataB <= 32'b00000100110010110010010000110100;
11'b00010010010: dataB <= 32'b01011111100011100110001111010010;
11'b00010010011: dataB <= 32'b00001010101100110110011010110111;
11'b00010010100: dataB <= 32'b00011110011000110011110101001011;
11'b00010010101: dataB <= 32'b00001000101001011000110000101100;
11'b00010010110: dataB <= 32'b01011001100010100110001111001111;
11'b00010010111: dataB <= 32'b00000010111000110000100101110111;
11'b00010011000: dataB <= 32'b01001101100010000110110101111100;
11'b00010011001: dataB <= 32'b00001000011110010011110101100101;
11'b00010011010: dataB <= 32'b11011110101101001111011110101010;
11'b00010011011: dataB <= 32'b00000101011101001111101101011011;
11'b00010011100: dataB <= 32'b11100111000101101010100100000011;
11'b00010011101: dataB <= 32'b00001000100010000100110101011101;
11'b00010011110: dataB <= 32'b01110011000001111111011101010100;
11'b00010011111: dataB <= 32'b00001000001000101000010001000111;
11'b00010100000: dataB <= 32'b10100111001001110001110100101010;
11'b00010100001: dataB <= 32'b00001101001100011001010011110100;
11'b00010100010: dataB <= 32'b11010011100110011010100111001101;
11'b00010100011: dataB <= 32'b00001000110001011011001111110010;
11'b00010100100: dataB <= 32'b10011111000001011111101001110100;
11'b00010100101: dataB <= 32'b00000100101001010110001110011011;
11'b00010100110: dataB <= 32'b11010101001001010101111011001101;
11'b00010100111: dataB <= 32'b00001010011010110011010001110011;
11'b00010101000: dataB <= 32'b00010000010110110100000110010101;
11'b00010101001: dataB <= 32'b00001111010101110010111101110001;
11'b00010101010: dataB <= 32'b01011111101111011110011011010100;
11'b00010101011: dataB <= 32'b00001011011101100111010110011110;
11'b00010101100: dataB <= 32'b10101001000011010100001010010110;
11'b00010101101: dataB <= 32'b00000101001001010110001001101111;
11'b00010101110: dataB <= 32'b00000011001001100100100100010111;
11'b00010101111: dataB <= 32'b00000000101111000110101100010100;
11'b00010110000: dataB <= 32'b10010011000111110100111100101110;
11'b00010110001: dataB <= 32'b00000001001010001100011101101011;
11'b00010110010: dataB <= 32'b01100011111001000101000001110111;
11'b00010110011: dataB <= 32'b00001010010001101110110010111111;
11'b00010110100: dataB <= 32'b11011100000101001101111010000101;
11'b00010110101: dataB <= 32'b00000101001111010110100101110000;
11'b00010110110: dataB <= 32'b10100001000010101101001000010111;
11'b00010110111: dataB <= 32'b00001000111110111010101110000101;
11'b00010111000: dataB <= 32'b01110010100100100101000011001111;
11'b00010111001: dataB <= 32'b00000100111011010111011011101010;
11'b00010111010: dataB <= 32'b10101010100011100011111110101000;
11'b00010111011: dataB <= 32'b00001001111110100111100010010011;
11'b00010111100: dataB <= 32'b11010010001011001110111001111101;
11'b00010111101: dataB <= 32'b00000011101110001010100000010101;
11'b00010111110: dataB <= 32'b01011111010010111011010110011001;
11'b00010111111: dataB <= 32'b00000011100100001010100001100110;
11'b00011000000: dataB <= 32'b01001110101111110100010111111011;
11'b00011000001: dataB <= 32'b00001100000011010111001100110100;
11'b00011000010: dataB <= 32'b11101100100101011101010110001111;
11'b00011000011: dataB <= 32'b00000010011000000011010001110110;
11'b00011000100: dataB <= 32'b10000010111101011001100010101111;
11'b00011000101: dataB <= 32'b00001101011010110011001100111011;
11'b00011000110: dataB <= 32'b00011010011111101101101010110100;
11'b00011000111: dataB <= 32'b00000011000100010110000101100011;
11'b00011001000: dataB <= 32'b01011101011011110011010111110011;
11'b00011001001: dataB <= 32'b00000011111001011100101110010100;
11'b00011001010: dataB <= 32'b00010101011011110100111100010100;
11'b00011001011: dataB <= 32'b00000101000110000011001010000011;
11'b00011001100: dataB <= 32'b10010011110111010010110110011101;
11'b00011001101: dataB <= 32'b00000111110111101100101110011011;
11'b00011001110: dataB <= 32'b11110010010001001100100111100001;
11'b00011001111: dataB <= 32'b00001001110111011111101001101101;
11'b00011010000: dataB <= 32'b11001000111011001100101101001101;
11'b00011010001: dataB <= 32'b00001000100100011010000101000011;
11'b00011010010: dataB <= 32'b01100000000101110111000111110111;
11'b00011010011: dataB <= 32'b00001100001101100101001101101001;
11'b00011010100: dataB <= 32'b10001001100000100100100001010101;
11'b00011010101: dataB <= 32'b00001000011110100101101101010011;
11'b00011010110: dataB <= 32'b10101011101101100100100111001110;
11'b00011010111: dataB <= 32'b00000110101001000010111110101111;
11'b00011011000: dataB <= 32'b00100110101000100110001000000001;
11'b00011011001: dataB <= 32'b00001010001010100000110111001001;
11'b00011011010: dataB <= 32'b10010001001101011100001000000101;
11'b00011011011: dataB <= 32'b00001011010100101110111100101110;
11'b00011011100: dataB <= 32'b11011011000010100101111001110001;
11'b00011011101: dataB <= 32'b00001111001101010011110101010110;
11'b00011011110: dataB <= 32'b10110000111101111011100011011001;
11'b00011011111: dataB <= 32'b00001000011000100101001110101111;
11'b00011100000: dataB <= 32'b10011110001001010010110011101111;
11'b00011100001: dataB <= 32'b00000000101110010000001100101100;
11'b00011100010: dataB <= 32'b10010011110110011110111010010110;
11'b00011100011: dataB <= 32'b00000100100111001010101110110010;
11'b00011100100: dataB <= 32'b00010101011010111000110011111001;
11'b00011100101: dataB <= 32'b00000000101100000011000110101010;
11'b00011100110: dataB <= 32'b10100000100001100011010001010101;
11'b00011100111: dataB <= 32'b00000101010100101000000100111101;
11'b00011101000: dataB <= 32'b01100111100011110100111111001101;
11'b00011101001: dataB <= 32'b00001001101010101110001111011110;
11'b00011101010: dataB <= 32'b00011000011100110100110100101101;
11'b00011101011: dataB <= 32'b00000111101001010110111000110101;
11'b00011101100: dataB <= 32'b01011111100110111101101110101001;
11'b00011101101: dataB <= 32'b00000100111011101010011010011111;
11'b00011101110: dataB <= 32'b10010101101110100110101000011101;
11'b00011101111: dataB <= 32'b00001011011101011101111001111101;
11'b00011110000: dataB <= 32'b00011010110001111111101101000101;
11'b00011110001: dataB <= 32'b00000111111110011001110101011100;
11'b00011110010: dataB <= 32'b00100111000001011010110010000110;
11'b00011110011: dataB <= 32'b00000110000010000101001001110110;
11'b00011110100: dataB <= 32'b10110010110010100111001101110000;
11'b00011110101: dataB <= 32'b00000110101000011110001101110111;
11'b00011110110: dataB <= 32'b01101001000001011010010100001101;
11'b00011110111: dataB <= 32'b00001100001000011101010111110011;
11'b00011111000: dataB <= 32'b10011011101110000010010110101110;
11'b00011111001: dataB <= 32'b00001001010000011111010011011001;
11'b00011111010: dataB <= 32'b01011111000010001111101010010011;
11'b00011111011: dataB <= 32'b00000011101100001100011010011011;
11'b00011111100: dataB <= 32'b00010111010001101110011010101011;
11'b00011111101: dataB <= 32'b00001100010111110101000001110100;
11'b00011111110: dataB <= 32'b10001010100010110011100111110110;
11'b00011111111: dataB <= 32'b00001111001111110000110001010001;
11'b00100000000: dataB <= 32'b11100111101011110101001011110001;
11'b00100000001: dataB <= 32'b00001101111001101011001110111101;
11'b00100000010: dataB <= 32'b10101000111011001011001011110100;
11'b00100000011: dataB <= 32'b00000100001100001100010110011111;
11'b00100000100: dataB <= 32'b01000111100001101100110110011001;
11'b00100000101: dataB <= 32'b00000000110101000101000000011101;
11'b00100000110: dataB <= 32'b11010111010011110011011100001010;
11'b00100000111: dataB <= 32'b00000000110000000110101101101011;
11'b00100001000: dataB <= 32'b01101111110101010101110011111011;
11'b00100001001: dataB <= 32'b00001010101111101010100111011110;
11'b00100001010: dataB <= 32'b00010000001001101110011000000100;
11'b00100001011: dataB <= 32'b00000101010001010010101101010001;
11'b00100001100: dataB <= 32'b01100001000010110100101001110110;
11'b00100001101: dataB <= 32'b00001011111101110100011010010101;
11'b00100001110: dataB <= 32'b00101100010100111110000011110011;
11'b00100001111: dataB <= 32'b00000111011100011101011111010001;
11'b00100010000: dataB <= 32'b01100010011111011010111100100100;
11'b00100010001: dataB <= 32'b00001100011011101011011010001011;
11'b00100010010: dataB <= 32'b11001010010111101101101100011010;
11'b00100010011: dataB <= 32'b00000011110010000110110100110110;
11'b00100010100: dataB <= 32'b10100011010010110010111000011010;
11'b00100010101: dataB <= 32'b00000010001000000110110110000110;
11'b00100010110: dataB <= 32'b00001100111111110010111001111010;
11'b00100010111: dataB <= 32'b00001001000001011011010000111101;
11'b00100011000: dataB <= 32'b11100110011101101101100110010001;
11'b00100011001: dataB <= 32'b00000100011011001001100110010110;
11'b00100011010: dataB <= 32'b10000101010101000010000011010100;
11'b00100011011: dataB <= 32'b00001110110101110100111100111100;
11'b00100011100: dataB <= 32'b10010100100011110100001011010010;
11'b00100011101: dataB <= 32'b00000001001000001100010001011011;
11'b00100011110: dataB <= 32'b00100001011011100001111000010011;
11'b00100011111: dataB <= 32'b00000101111100011000110010010100;
11'b00100100000: dataB <= 32'b00011011100011110011011100110000;
11'b00100100001: dataB <= 32'b00000011101001000111100001111011;
11'b00100100010: dataB <= 32'b01011111111010111001111001011101;
11'b00100100011: dataB <= 32'b00001001010110101000100010010011;
11'b00100100100: dataB <= 32'b00100110000101010101010100100010;
11'b00100100101: dataB <= 32'b00001011010101101001100110000110;
11'b00100100110: dataB <= 32'b10001001001011001011101100001001;
11'b00100100111: dataB <= 32'b00000110100101010000001101001100;
11'b00100101000: dataB <= 32'b11010100001010011110111001010110;
11'b00100101001: dataB <= 32'b00001011101010100111001001001001;
11'b00100101010: dataB <= 32'b00010001101100110101100010111010;
11'b00100101011: dataB <= 32'b00001010111101101101100101010100;
11'b00100101100: dataB <= 32'b11110011100001110100110111001110;
11'b00100101101: dataB <= 32'b00000101001010000011010111010110;
11'b00100101110: dataB <= 32'b01100010100101000110110101000001;
11'b00100101111: dataB <= 32'b00001001001001011110110110100000;
11'b00100110000: dataB <= 32'b01010101011001100100100110000110;
11'b00100110001: dataB <= 32'b00001011110001101100110001010111;
11'b00100110010: dataB <= 32'b01011011000110111101011010001111;
11'b00100110011: dataB <= 32'b00001110000111011111111001111111;
11'b00100110100: dataB <= 32'b11101110110001111011100101011100;
11'b00100110101: dataB <= 32'b00001001110111100111001011010110;
11'b00100110110: dataB <= 32'b10010100001101001011010100010010;
11'b00100110111: dataB <= 32'b00000000110100001000011100111101;
11'b00100111000: dataB <= 32'b00011111111010111110011011110100;
11'b00100111001: dataB <= 32'b00000011001011001000111110011010;
11'b00100111010: dataB <= 32'b11011011011110001000010101111100;
11'b00100111011: dataB <= 32'b00000000110001000101011110001001;
11'b00100111100: dataB <= 32'b01011010100101100011110010111010;
11'b00100111101: dataB <= 32'b00000110010110011110000101011110;
11'b00100111110: dataB <= 32'b00101011011011110011011110000111;
11'b00100111111: dataB <= 32'b00001000101001100010000111110101;
11'b00101000000: dataB <= 32'b11010010100101000101100100010000;
11'b00101000001: dataB <= 32'b00000110101010010101000001000101;
11'b00101000010: dataB <= 32'b10100111100011001100101101000100;
11'b00101000011: dataB <= 32'b00000111011100100010010111000110;
11'b00101000100: dataB <= 32'b10011111110111000101111010111100;
11'b00101000101: dataB <= 32'b00001101111010101001111010001101;
11'b00101000110: dataB <= 32'b10011000110110101111101010100010;
11'b00101000111: dataB <= 32'b00001010111101100101110101100100;
11'b00101001000: dataB <= 32'b00100110111001010011010000101100;
11'b00101001001: dataB <= 32'b00000011100101001001011110010110;
11'b00101001010: dataB <= 32'b10101110100111001110011101001100;
11'b00101001011: dataB <= 32'b00000101101001010110010010100111;
11'b00101001100: dataB <= 32'b11101000111001000010110011110000;
11'b00101001101: dataB <= 32'b00001010100101100001010111100001;
11'b00101001110: dataB <= 32'b10100011101101110010010110101111;
11'b00101001111: dataB <= 32'b00001001001111100011010010110000;
11'b00101010000: dataB <= 32'b00011111000010111111011010110001;
11'b00101010001: dataB <= 32'b00000011010000000110101010001011;
11'b00101010010: dataB <= 32'b00011011010110001110011001101001;
11'b00101010011: dataB <= 32'b00001101010100110010110001110100;
11'b00101010100: dataB <= 32'b01000110110110100010111000110110;
11'b00101010101: dataB <= 32'b00001110101001101100100100111010;
11'b00101010110: dataB <= 32'b11101111100011110011111011101110;
11'b00101010111: dataB <= 32'b00001111010100101101000111001100;
11'b00101011000: dataB <= 32'b00011100101101100001101010001000;
11'b00101011001: dataB <= 32'b00000110010111001011100111110011;
11'b00101011010: dataB <= 32'b00110001110010011100101100110011;
11'b00101011011: dataB <= 32'b00001010111110100001110110101111;
11'b00101011100: dataB <= 32'b10101001010001101000010101000111;
11'b00101011101: dataB <= 32'b00001000011110010111110001111100;
11'b00101011110: dataB <= 32'b00111010100010111101011101111000;
11'b00101011111: dataB <= 32'b00000111101010010010101011001001;
11'b00101100000: dataB <= 32'b01000101011111001100100010001111;
11'b00101100001: dataB <= 32'b00001000110101010111011000100101;
11'b00101100010: dataB <= 32'b01100000111110010010011011001100;
11'b00101100011: dataB <= 32'b00001110101000001100010110101011;
11'b00101100100: dataB <= 32'b01001010100111000110001001111000;
11'b00101100101: dataB <= 32'b00001110010001101111000100100001;
11'b00101100110: dataB <= 32'b10001110111001011001000010000110;
11'b00101100111: dataB <= 32'b00001101100111101100101001101011;
11'b00101101000: dataB <= 32'b01001011101010110000101101000111;
11'b00101101001: dataB <= 32'b00001001011000011011110011011110;
11'b00101101010: dataB <= 32'b11101000111001011010011101001111;
11'b00101101011: dataB <= 32'b00000100011011011011110011010011;
11'b00101101100: dataB <= 32'b00011111100101011000011101001100;
11'b00101101101: dataB <= 32'b00000000101101101001001010100110;
11'b00101101110: dataB <= 32'b01001110110010110100101000110011;
11'b00101101111: dataB <= 32'b00001101110111110011101111011011;
11'b00101110000: dataB <= 32'b00101011110101000101111010011001;
11'b00101110001: dataB <= 32'b00001010100010011110010110010110;
11'b00101110010: dataB <= 32'b00010001010110000000011001001001;
11'b00101110011: dataB <= 32'b00000100011101001001100101110101;
11'b00101110100: dataB <= 32'b01101100111100111000111001101111;
11'b00101110101: dataB <= 32'b00001110010100011001001110000011;
11'b00101110110: dataB <= 32'b00110001001001101000011000000110;
11'b00101110111: dataB <= 32'b00000100111000110001110001100100;
11'b00101111000: dataB <= 32'b01111101000000111010001110101101;
11'b00101111001: dataB <= 32'b00001011001101010000101101101011;
11'b00101111010: dataB <= 32'b11000010110010101101010001010110;
11'b00101111011: dataB <= 32'b00001010101001110010101111000011;
11'b00101111100: dataB <= 32'b10100101101101110001100100100111;
11'b00101111101: dataB <= 32'b00000010110010000111011110010101;
11'b00101111110: dataB <= 32'b10000101010111011011001011001101;
11'b00101111111: dataB <= 32'b00000101001000100100110000111101;
11'b00110000000: dataB <= 32'b01110111011110110110011101011010;
11'b00110000001: dataB <= 32'b00001110101010110010100110000101;
11'b00110000010: dataB <= 32'b01110000011010011100010111010001;
11'b00110000011: dataB <= 32'b00000101010101101011111011011001;
11'b00110000100: dataB <= 32'b11010010111011011101110000110101;
11'b00110000101: dataB <= 32'b00000100101101011011000000001010;
11'b00110000110: dataB <= 32'b01101101010110010100110011010011;
11'b00110000111: dataB <= 32'b00001000101000011000100111101101;
11'b00110001000: dataB <= 32'b00100011001010101010000111101011;
11'b00110001001: dataB <= 32'b00000011100011111101000011101100;
11'b00110001010: dataB <= 32'b01011000100001110100001110010101;
11'b00110001011: dataB <= 32'b00001011101100100100110011011001;
11'b00110001100: dataB <= 32'b00000111010101101101101001010111;
11'b00110001101: dataB <= 32'b00001010011110001111101110110110;
11'b00110001110: dataB <= 32'b00111101000011001010001010001000;
11'b00110001111: dataB <= 32'b00000101111001011111101101000011;
11'b00110010000: dataB <= 32'b10101111001000001011101110010100;
11'b00110010001: dataB <= 32'b00001000111110101111110100111011;
11'b00110010010: dataB <= 32'b00010011001001111100111101011010;
11'b00110010011: dataB <= 32'b00001011010011000011000011001101;
11'b00110010100: dataB <= 32'b01101100101001101000010011100011;
11'b00110010101: dataB <= 32'b00000100101110000010111010100000;
11'b00110010110: dataB <= 32'b11010011011010110101111000010111;
11'b00110010111: dataB <= 32'b00000101010010100001010110111101;
11'b00110011000: dataB <= 32'b11110000110010010001100010000101;
11'b00110011001: dataB <= 32'b00001110010001001010111011010001;
11'b00110011010: dataB <= 32'b10111011000010111001111110001010;
11'b00110011011: dataB <= 32'b00001101000100111100101110110011;
11'b00110011100: dataB <= 32'b11011011001111110010100001001010;
11'b00110011101: dataB <= 32'b00001110101010111010110110010100;
11'b00110011110: dataB <= 32'b01011100110001101101010110011110;
11'b00110011111: dataB <= 32'b00000010111000101111101111000011;
11'b00110100000: dataB <= 32'b11010010100011001001100110000101;
11'b00110100001: dataB <= 32'b00000100110100001001010011110010;
11'b00110100010: dataB <= 32'b11011100101101011101111000011000;
11'b00110100011: dataB <= 32'b00000010101010101010111100111000;
11'b00110100100: dataB <= 32'b01110110111001001100010111110010;
11'b00110100101: dataB <= 32'b00000111101101101000111000010010;
11'b00110100110: dataB <= 32'b10100001000011101010001000101010;
11'b00110100111: dataB <= 32'b00001000011001010101110001100011;
11'b00110101000: dataB <= 32'b01101011001011001011100100101100;
11'b00110101001: dataB <= 32'b00001010000101011000011010000100;
11'b00110101010: dataB <= 32'b00011011110001011010111011001110;
11'b00110101011: dataB <= 32'b00000100100010010010100101001110;
11'b00110101100: dataB <= 32'b10110000100001111000010111001000;
11'b00110101101: dataB <= 32'b00001010000001100010100110011001;
11'b00110101110: dataB <= 32'b10100000101110000001011011001011;
11'b00110101111: dataB <= 32'b00000100110101000101010011110100;
11'b00110110000: dataB <= 32'b01100101111010010100111011110111;
11'b00110110001: dataB <= 32'b00000111111110010111110010000111;
11'b00110110010: dataB <= 32'b10100011011010011000010111000110;
11'b00110110011: dataB <= 32'b00000101011101001111100101110100;
11'b00110110100: dataB <= 32'b00111100111010100101111011111100;
11'b00110110101: dataB <= 32'b00001000101011011000100011101010;
11'b00110110110: dataB <= 32'b01000011000110111101100010101011;
11'b00110110111: dataB <= 32'b00000111110101010011010000011100;
11'b00110111000: dataB <= 32'b11100000111110100010101011101111;
11'b00110111001: dataB <= 32'b00001111001110010110001010110011;
11'b00110111010: dataB <= 32'b10010010011010100110110111111001;
11'b00110111011: dataB <= 32'b00001101110110101101010001001000;
11'b00110111100: dataB <= 32'b01010000101001111000110100000010;
11'b00110111101: dataB <= 32'b00001111001100110000110001110011;
11'b00110111110: dataB <= 32'b01000101011011011001101110101100;
11'b00110111111: dataB <= 32'b00000111011000010001101010111111;
11'b00111000000: dataB <= 32'b11101001000001101010001100110011;
11'b00111000001: dataB <= 32'b00000010011000010001101011001100;
11'b00111000010: dataB <= 32'b01010111100010001000011101110000;
11'b00111000011: dataB <= 32'b00000001100111100111010010001110;
11'b00111000100: dataB <= 32'b01010010100110101101000111110011;
11'b00111000101: dataB <= 32'b00001100011011101001111011011100;
11'b00111000110: dataB <= 32'b00011111111000110101000111111010;
11'b00111000111: dataB <= 32'b00001101000101100110011001110110;
11'b00111001000: dataB <= 32'b11001111001010110000101010001010;
11'b00111001001: dataB <= 32'b00000010011001000011010001100100;
11'b00111001010: dataB <= 32'b01101101000101101000011001110000;
11'b00111001011: dataB <= 32'b00001100111000010111000110001011;
11'b00111001100: dataB <= 32'b11101101010110011000011010000111;
11'b00111001101: dataB <= 32'b00000011010101100101111001100011;
11'b00111001110: dataB <= 32'b00111011011001011001011110110011;
11'b00111001111: dataB <= 32'b00001011110000010110100101110011;
11'b00111010000: dataB <= 32'b10001000011010010101100000110000;
11'b00111010001: dataB <= 32'b00001011101100110101000010111100;
11'b00111010010: dataB <= 32'b11011101101110010001100110100101;
11'b00111010011: dataB <= 32'b00000010001110000011001001111101;
11'b00111010100: dataB <= 32'b10000010111111100100011011110000;
11'b00111010101: dataB <= 32'b00000110100111100110110100101100;
11'b00111010110: dataB <= 32'b01110001101110010110111010111101;
11'b00111010111: dataB <= 32'b00001111001111110110110101110101;
11'b00111011000: dataB <= 32'b10110110101010010100110111010001;
11'b00111011001: dataB <= 32'b00000100110010011111111011110010;
11'b00111011010: dataB <= 32'b10010100110011000110110000101111;
11'b00111011011: dataB <= 32'b00000101001011011010111100100001;
11'b00111011100: dataB <= 32'b10100111011110000101000010101111;
11'b00111011101: dataB <= 32'b00001010001001011110100011010110;
11'b00111011110: dataB <= 32'b01100001001010111010111000101100;
11'b00111011111: dataB <= 32'b00000110100001111011011011011101;
11'b00111100000: dataB <= 32'b10011110011101110100001100111001;
11'b00111100001: dataB <= 32'b00001100001111100110110111110010;
11'b00111100010: dataB <= 32'b10000101000001011101010111111000;
11'b00111100011: dataB <= 32'b00000111011110000111011110010110;
11'b00111100100: dataB <= 32'b01111011011011011011001011001011;
11'b00111100101: dataB <= 32'b00000011110110010111101001010010;
11'b00111100110: dataB <= 32'b10101101010100011010001100111000;
11'b00111100111: dataB <= 32'b00000110011110100011111001000010;
11'b00111101000: dataB <= 32'b00010000111101101100111010111101;
11'b00111101001: dataB <= 32'b00001010010101000010101110110110;
11'b00111101010: dataB <= 32'b00110000110010011000010110100001;
11'b00111101011: dataB <= 32'b00000101001100000110100011001001;
11'b00111101100: dataB <= 32'b01001111001110011110010110110110;
11'b00111101101: dataB <= 32'b00000100110000011101010010100110;
11'b00111101110: dataB <= 32'b00110011000010110010000100100010;
11'b00111101111: dataB <= 32'b00001101110110001100101011101011;
11'b00111110000: dataB <= 32'b00110111010111010010111110101111;
11'b00111110001: dataB <= 32'b00001110101001111101000110110100;
11'b00111110010: dataB <= 32'b00011001001011110100000010100101;
11'b00111110011: dataB <= 32'b00001111010000111011001110000101;
11'b00111110100: dataB <= 32'b01100000110001011101000011011011;
11'b00111110101: dataB <= 32'b00000001010011100101110111000100;
11'b00111110110: dataB <= 32'b01011000011011100010111000000100;
11'b00111110111: dataB <= 32'b00000100010010000111000011110100;
11'b00111111000: dataB <= 32'b01100000101101001101000110110111;
11'b00111111001: dataB <= 32'b00000100000111101011000101101000;
11'b00111111010: dataB <= 32'b00110111001001001011110111010010;
11'b00111111011: dataB <= 32'b00001000001101101001000000110001;
11'b00111111100: dataB <= 32'b00100001000011110011101001101011;
11'b00111111101: dataB <= 32'b00000110011000001101100101101011;
11'b00111111110: dataB <= 32'b01101001010011001100100101101010;
11'b00111111111: dataB <= 32'b00001011100111100000010110000100;
11'b01000000000: dataB <= 32'b01010001101001110010011011010000;
11'b01000000001: dataB <= 32'b00000111100001011000011100110101;
11'b01000000010: dataB <= 32'b00110100110010100000011000101000;
11'b01000000011: dataB <= 32'b00001100100100100110101010111010;
11'b01000000100: dataB <= 32'b11100100110010100001101100001110;
11'b01000000101: dataB <= 32'b00000100010010000010111011100101;
11'b01000000110: dataB <= 32'b00011011111010000101001001111001;
11'b01000000111: dataB <= 32'b00000100111101001101100101011111;
11'b01000001000: dataB <= 32'b01011111011011000000111000100110;
11'b01000001001: dataB <= 32'b00000010111010001001010101101100;
11'b01000001010: dataB <= 32'b10111101010010001110001001011110;
11'b01000001011: dataB <= 32'b00001001101100011110011111110011;
11'b01000001100: dataB <= 32'b00000010110010100110000100000111;
11'b01000001101: dataB <= 32'b00000110110101010001000100011011;
11'b01000001110: dataB <= 32'b01100000111110110011001011110010;
11'b01000001111: dataB <= 32'b00001111010100100010000110110100;
11'b01000010000: dataB <= 32'b01011010010001111111000110011000;
11'b01000010001: dataB <= 32'b00001100011010101001011001111000;
11'b01000010010: dataB <= 32'b00010100100010100001000111000001;
11'b01000010011: dataB <= 32'b00001111010010110001000001111011;
11'b01000010100: dataB <= 32'b10000011000011110010111110110001;
11'b01000010101: dataB <= 32'b00000101110111001011011110001111;
11'b01000010110: dataB <= 32'b10100111001010000010001100010110;
11'b01000010111: dataB <= 32'b00000001010011001011011111000101;
11'b01000011000: dataB <= 32'b00010011010110111000101101010100;
11'b01000011001: dataB <= 32'b00000011100011100011010101101110;
11'b01000011010: dataB <= 32'b10011000011110011101100111010011;
11'b01000011011: dataB <= 32'b00001001111101011101111011010101;
11'b01000011100: dataB <= 32'b11010101110100101100000101111001;
11'b01000011101: dataB <= 32'b00001110101010101110100001011101;
11'b01000011110: dataB <= 32'b01001100111011011001101011001100;
11'b01000011111: dataB <= 32'b00000000110011000010111001011100;
11'b01000100000: dataB <= 32'b10101001001110010000011001010001;
11'b01000100001: dataB <= 32'b00001010111011010110111110010011;
11'b01000100010: dataB <= 32'b10101001100011000000111011001010;
11'b01000100011: dataB <= 32'b00000010010001011011111001101011;
11'b01000100100: dataB <= 32'b00110011101101111001001101111000;
11'b01000100101: dataB <= 32'b00001011010010011100011101111011;
11'b01000100110: dataB <= 32'b01010000001110000101110000101010;
11'b01000100111: dataB <= 32'b00001100001111110011010010110101;
11'b01000101000: dataB <= 32'b10010011101010101010001000100101;
11'b01000101001: dataB <= 32'b00000011001010000010110001101101;
11'b01000101010: dataB <= 32'b10000100101011011101011011010010;
11'b01000101011: dataB <= 32'b00001000100110101000111100101011;
11'b01000101100: dataB <= 32'b00100111110101101110110111111110;
11'b01000101101: dataB <= 32'b00001110110101110111001001100101;
11'b01000101110: dataB <= 32'b00111000111010001100110110110000;
11'b01000101111: dataB <= 32'b00000100010000010011110111110100;
11'b01000110000: dataB <= 32'b10011000101010011111010001001001;
11'b01000110001: dataB <= 32'b00000110001001011100111001001000;
11'b01000110010: dataB <= 32'b01100001100001111101000011001011;
11'b01000110011: dataB <= 32'b00001011001011100100100010101111;
11'b01000110100: dataB <= 32'b01011111001011000011101001001100;
11'b01000110101: dataB <= 32'b00001001000001110011101111000110;
11'b01000110110: dataB <= 32'b00100110011101110011111010011100;
11'b01000110111: dataB <= 32'b00001100010011101000111111110100;
11'b01000111000: dataB <= 32'b10000110101101001100110110010111;
11'b01000111001: dataB <= 32'b00000100011101000011001001110110;
11'b01000111010: dataB <= 32'b00110011101111011100011100001110;
11'b01000111011: dataB <= 32'b00000011010011001111011101101010;
11'b01000111100: dataB <= 32'b00100111011100110001001010111011;
11'b01000111101: dataB <= 32'b00000011011011010111111001010010;
11'b01000111110: dataB <= 32'b01010010110101100100100111111110;
11'b01000111111: dataB <= 32'b00001001010110001000011010011110;
11'b01001000000: dataB <= 32'b01110001000011000000111001000001;
11'b01001000001: dataB <= 32'b00000110001010001100010011101010;
11'b01001000010: dataB <= 32'b10001101000001111110010101110101;
11'b01001000011: dataB <= 32'b00000100101110011001001110000110;
11'b01001000100: dataB <= 32'b01110001001111000010110111100001;
11'b01001000101: dataB <= 32'b00001100011010010010011111101100;
11'b01001000110: dataB <= 32'b11110001100111011011111110010100;
11'b01001000111: dataB <= 32'b00001111001111111011011010101100;
11'b01001001000: dataB <= 32'b00010111000011101101100101000010;
11'b01001001001: dataB <= 32'b00001110110101110111100001111101;
11'b01001001010: dataB <= 32'b00100010110001010100100001110111;
11'b01001001011: dataB <= 32'b00000001001110011011110110111101;
11'b01001001100: dataB <= 32'b11100000011011101100001010000101;
11'b01001001101: dataB <= 32'b00000100001111001000101111101101;
11'b01001001110: dataB <= 32'b01100100110000111100010101010110;
11'b01001001111: dataB <= 32'b00000110000101101001001110010000;
11'b01001010000: dataB <= 32'b01110011011001010011000110110001;
11'b01001010001: dataB <= 32'b00001000101110100111001001011000;
11'b01001010010: dataB <= 32'b00100001000011110101001010001100;
11'b01001010011: dataB <= 32'b00000100110110000111010001110011;
11'b01001010100: dataB <= 32'b01100101010110111101010110101001;
11'b01001010101: dataB <= 32'b00001101001011101000011001111100;
11'b01001010110: dataB <= 32'b01001011011110000010011010110011;
11'b01001010111: dataB <= 32'b00001010100001011110011000100100;
11'b01001011000: dataB <= 32'b00110111000011001001001010001001;
11'b01001011001: dataB <= 32'b00001110101001101010110011001011;
11'b01001011010: dataB <= 32'b00100110110110111010011100010001;
11'b01001011011: dataB <= 32'b00000011101111000110100111000111;
11'b01001011100: dataB <= 32'b01001111110001110101000111111010;
11'b01001011101: dataB <= 32'b00000010011010000111010100110110;
11'b01001011110: dataB <= 32'b00011011010111100001111010100111;
11'b01001011111: dataB <= 32'b00000001010101000101000001101100;
11'b01001100000: dataB <= 32'b00110111100101101110000110011101;
11'b01001100001: dataB <= 32'b00001010001110100100100011110101;
11'b01001100010: dataB <= 32'b11001000011010000110100101100101;
11'b01001100011: dataB <= 32'b00000101110011010000111000110001;
11'b01001100100: dataB <= 32'b00100000111110111011111011010100;
11'b01001100101: dataB <= 32'b00001101111001101100001110100101;
11'b01001100110: dataB <= 32'b01100010010001011110110100110110;
11'b01001100111: dataB <= 32'b00001001111100100011011110101000;
11'b01001101000: dataB <= 32'b00011100011111000001111010000001;
11'b01001101001: dataB <= 32'b00001110010111101111001110000011;
11'b01001101010: dataB <= 32'b10000010101011110100001101110110;
11'b01001101011: dataB <= 32'b00000100010101000111001001011111;
11'b01001101100: dataB <= 32'b01100101001110011010011010011001;
11'b01001101101: dataB <= 32'b00000001001101000111001010100110;
11'b01001101110: dataB <= 32'b11001111001011011001101011111000;
11'b01001101111: dataB <= 32'b00000110100001011111010101010101;
11'b01001110000: dataB <= 32'b01100000011010000101110110110010;
11'b01001110001: dataB <= 32'b00000110111101010001110110111110;
11'b01001110010: dataB <= 32'b01001011101000110010110100010111;
11'b01001110011: dataB <= 32'b00001111010000110010110001000101;
11'b01001110100: dataB <= 32'b11001110101111110010111011101111;
11'b01001110101: dataB <= 32'b00000000101110000100100001010011;
11'b01001110110: dataB <= 32'b11100111010111000000111000110010;
11'b01001110111: dataB <= 32'b00001000011101010110110110010011;
11'b01001111000: dataB <= 32'b01100001100111100001111100001101;
11'b01001111001: dataB <= 32'b00000010101101001111110001110011;
11'b01001111010: dataB <= 32'b00101001111010011001011011111011;
11'b01001111011: dataB <= 32'b00001010110101100010011110001011;
11'b01001111100: dataB <= 32'b11011100000101101101100010000101;
11'b01001111101: dataB <= 32'b00001011110010101111011110011101;
11'b01001111110: dataB <= 32'b01001101011111000010111010100110;
11'b01001111111: dataB <= 32'b00000100100111001000011101010101;
11'b01010000000: dataB <= 32'b10001010010111000110011010110101;
11'b01010000001: dataB <= 32'b00001010000111101001000100110010;
11'b01010000010: dataB <= 32'b10011011110101001110010101011101;
11'b01010000011: dataB <= 32'b00001101011010110011011001011100;
11'b01010000100: dataB <= 32'b10110111001101111101000110101111;
11'b01010000101: dataB <= 32'b00000100101101001001101011101101;
11'b01010000110: dataB <= 32'b01011100100101101111010010100100;
11'b01010000111: dataB <= 32'b00000111101000011100111001111000;
11'b01010001000: dataB <= 32'b10011011011101101100110100101000;
11'b01010001001: dataB <= 32'b00001011101110101000100101111111;
11'b01010001010: dataB <= 32'b00011101001011000100101001101110;
11'b01010001011: dataB <= 32'b00001100000011101001111010100111;
11'b01010001100: dataB <= 32'b10101010100101110011110111111101;
11'b01010001101: dataB <= 32'b00001011010101101001000111101101;
11'b01010001110: dataB <= 32'b01001100011001000100000100110101;
11'b01010001111: dataB <= 32'b00000010011001000100110001010110;
11'b01010010000: dataB <= 32'b11101001111011010101101100010001;
11'b01010010001: dataB <= 32'b00000010101111001011010010000001;
11'b01010010010: dataB <= 32'b11100001100001100000011000011101;
11'b01010010011: dataB <= 32'b00000001010111001101101101110001;
11'b01010010100: dataB <= 32'b10010100101001100100000101011101;
11'b01010010101: dataB <= 32'b00000111110111010010001001111110;
11'b01010010110: dataB <= 32'b11101111001111100001111100000011;
11'b01010010111: dataB <= 32'b00000111001001011000000111110011;
11'b01010011000: dataB <= 32'b01001110110001011110010100110011;
11'b01010011001: dataB <= 32'b00000101101011010111000101011110;
11'b01010011010: dataB <= 32'b10101101011011010011111010100001;
11'b01010011011: dataB <= 32'b00001001111100011000010111011101;
11'b01010011100: dataB <= 32'b01101001110011010100111100111001;
11'b01010011101: dataB <= 32'b00001111010101110011101110100101;
11'b01010011110: dataB <= 32'b11010110111011010110101000000001;
11'b01010011111: dataB <= 32'b00001101011010101111101101101100;
11'b01010100000: dataB <= 32'b11100100110101001100000000110001;
11'b01010100001: dataB <= 32'b00000010001001010001101110101101;
11'b01010100010: dataB <= 32'b11101000011011100101011100001000;
11'b01010100011: dataB <= 32'b00000100101100001110011111001110;
11'b01010100100: dataB <= 32'b11100110110100111011100100010011;
11'b01010100101: dataB <= 32'b00001000000100100101010011000000;
11'b01010100110: dataB <= 32'b01101101101001011010100110110000;
11'b01010100111: dataB <= 32'b00001000101110100101001110000000;
11'b01010101000: dataB <= 32'b11100001000011011110011010101110;
11'b01010101001: dataB <= 32'b00000011110011000100111110000010;
11'b01010101010: dataB <= 32'b01100001011010100110001000001000;
11'b01010101011: dataB <= 32'b00001101101111101110100101111100;
11'b01010101100: dataB <= 32'b01000111001010010010101010010101;
11'b01010101101: dataB <= 32'b00001101000100100110011100101011;
11'b01010101110: dataB <= 32'b00110101010111101010011011001011;
11'b01010101111: dataB <= 32'b00001111001111101100111011010100;
11'b01010110000: dataB <= 32'b11011010110001001010001000100111;
11'b01010110001: dataB <= 32'b00000111111000010011110011100001;
11'b01010110010: dataB <= 32'b01111001100010100100011101010000;
11'b01010110011: dataB <= 32'b00001101011011101011110011001110;
11'b01010110100: dataB <= 32'b10101011001000111000110011101010;
11'b01010110101: dataB <= 32'b00001010111101100001110110000100;
11'b01010110110: dataB <= 32'b01110010010011000100101110110011;
11'b01010110111: dataB <= 32'b00000111001011010000110110100000;
11'b01010111000: dataB <= 32'b01001101101111010011110010110100;
11'b01010111001: dataB <= 32'b00001001110100011101011100111110;
11'b01010111010: dataB <= 32'b11011110111101111010001010001001;
11'b01010111011: dataB <= 32'b00001100100100000110100110100010;
11'b01010111100: dataB <= 32'b10001000111011011101001011010110;
11'b01010111101: dataB <= 32'b00001110001100101110111000001010;
11'b01010111110: dataB <= 32'b11001111000100111001110000101011;
11'b01010111111: dataB <= 32'b00001011100011100110100001100011;
11'b01011000000: dataB <= 32'b00010101111010000000011011000100;
11'b01011000001: dataB <= 32'b00001010110111100101110011110101;
11'b01011000010: dataB <= 32'b11100110110101001011001100101011;
11'b01011000011: dataB <= 32'b00000110111101100101110011001010;
11'b01011000100: dataB <= 32'b01100101100000110001001100001000;
11'b01011000101: dataB <= 32'b00000000110010101011000010111101;
11'b01011000110: dataB <= 32'b00001100111110111011111001010010;
11'b01011000111: dataB <= 32'b00001110110010111011011111001010;
11'b01011001000: dataB <= 32'b11110101101001011110011011110111;
11'b01011001001: dataB <= 32'b00001000000001011000011010101101;
11'b01011001010: dataB <= 32'b01010111100001011000010111101000;
11'b01011001011: dataB <= 32'b00000111011110010001110101111101;
11'b01011001100: dataB <= 32'b01101010110000011001111001001110;
11'b01011001101: dataB <= 32'b00001110101111011011010001111011;
11'b01011001110: dataB <= 32'b01110010111100111000110110100111;
11'b01011001111: dataB <= 32'b00000110111010111001100001101100;
11'b01011010000: dataB <= 32'b10111100101100101011001101101000;
11'b01011010001: dataB <= 32'b00001010101010001110111001100011;
11'b01011010010: dataB <= 32'b00000011000110110100100010111011;
11'b01011010011: dataB <= 32'b00001001001000101110100010111011;
11'b01011010100: dataB <= 32'b01101111100101011001110011001010;
11'b01011010101: dataB <= 32'b00000011110110001111101110101101;
11'b01011010110: dataB <= 32'b01001011101011001001111010101010;
11'b01011010111: dataB <= 32'b00000011101011100010101101010110;
11'b01011011000: dataB <= 32'b00111011001011001101101110110101;
11'b01011011001: dataB <= 32'b00001101000101101100011010010101;
11'b01011011010: dataB <= 32'b10100110010010100100000111110010;
11'b01011011011: dataB <= 32'b00000110110110110101101110110000;
11'b01011011100: dataB <= 32'b00010011000111101100100010011010;
11'b01011011101: dataB <= 32'b00000100010000011101000100001100;
11'b01011011110: dataB <= 32'b00101111001010011100100100010110;
11'b01011011111: dataB <= 32'b00000111001000010010101111110100;
11'b01011100000: dataB <= 32'b11100101000110010001110111001100;
11'b01011100001: dataB <= 32'b00000001100111111100101111100010;
11'b01011100010: dataB <= 32'b10010010101001111100011110110000;
11'b01011100011: dataB <= 32'b00001010101001100010101110110000;
11'b01011100100: dataB <= 32'b01001101100110000101111010110110;
11'b01011100101: dataB <= 32'b00001100111011011001110111001101;
11'b01011100110: dataB <= 32'b11111100101110110001011000100111;
11'b01011100111: dataB <= 32'b00000111111010101001101000111011;
11'b01011101000: dataB <= 32'b01110000111100001100111110101111;
11'b01011101001: dataB <= 32'b00001011111101110111100100111100;
11'b01011101010: dataB <= 32'b00010101010110000100111110110101;
11'b01011101011: dataB <= 32'b00001011110000000101011011010100;
11'b01011101100: dataB <= 32'b01100110100000111000110001100111;
11'b01011101101: dataB <= 32'b00000100110001000011001101111000;
11'b01011101110: dataB <= 32'b00011001100011001101001001110110;
11'b01011101111: dataB <= 32'b00000101110100100011010011001101;
11'b01011110000: dataB <= 32'b00101100100101111001010000101010;
11'b01011110001: dataB <= 32'b00001110001100001011001110110001;
11'b01011110010: dataB <= 32'b11111000101110011001011100100110;
11'b01011110011: dataB <= 32'b00001010100001110110011010101010;
11'b01011110100: dataB <= 32'b10011101010011010001010000101111;
11'b01011110101: dataB <= 32'b00001101000101110110100010011100;
11'b01011110110: dataB <= 32'b10011010110110000101101000111110;
11'b01011110111: dataB <= 32'b00000100111011110111011110111010;
11'b01011111000: dataB <= 32'b10001100101110101000110100000111;
11'b01011111001: dataB <= 32'b00000110010110001111100011011001;
11'b01011111010: dataB <= 32'b11011010110001110110001001110111;
11'b01011111011: dataB <= 32'b00000010001111101000110100011001;
11'b01011111100: dataB <= 32'b11110100100101010101001000010010;
11'b01011111101: dataB <= 32'b00000111001110100110110100001011;
11'b01011111110: dataB <= 32'b11100000111111001001000111001010;
11'b01011111111: dataB <= 32'b00001001111000011111110101011011;
11'b01100000000: dataB <= 32'b00101100111111000010110100001111;
11'b01100000001: dataB <= 32'b00000111100100010010100010001100;
11'b01100000010: dataB <= 32'b10100101110001010011011010101011;
11'b01100000011: dataB <= 32'b00000010000101001110110001101110;
11'b01100000100: dataB <= 32'b01101010010101001000100101101001;
11'b01100000101: dataB <= 32'b00000111100001011100100110000001;
11'b01100000110: dataB <= 32'b11011000110100110010110111000111;
11'b01100000111: dataB <= 32'b00001001010111011101111010111000;
11'b01100001000: dataB <= 32'b00111101001010100011111100101100;
11'b01100001001: dataB <= 32'b00001110110110110011100111100101;
11'b01100001010: dataB <= 32'b10101101000000011001110011001110;
11'b01100001011: dataB <= 32'b00001101011010101011101110001100;
11'b01100001100: dataB <= 32'b01101000000111000011101111001101;
11'b01100001101: dataB <= 32'b00000110001100001111000001110000;
11'b01100001110: dataB <= 32'b00011001111011000010110011110111;
11'b01100001111: dataB <= 32'b00001010110010100011011101100111;
11'b01100010000: dataB <= 32'b01011110111101100010011001001000;
11'b01100010001: dataB <= 32'b00001010000001000010111010001010;
11'b01100010010: dataB <= 32'b00001001001011100100001100010011;
11'b01100010011: dataB <= 32'b00001101000111101100101100001100;
11'b01100010100: dataB <= 32'b00010001010100100010110000110001;
11'b01100010101: dataB <= 32'b00001001000001100000011101100100;
11'b01100010110: dataB <= 32'b10100001111001011000011000100010;
11'b01100010111: dataB <= 32'b00001011110100101111101011110011;
11'b01100011000: dataB <= 32'b11100100110001000011111011000111;
11'b01100011001: dataB <= 32'b00001001111101101111101010110001;
11'b01100011010: dataB <= 32'b10101011011000010010001010000101;
11'b01100011011: dataB <= 32'b00000001111000101010111011000100;
11'b01100011100: dataB <= 32'b01001111001110110011001001110001;
11'b01100011101: dataB <= 32'b00001110101100111101000110110001;
11'b01100011110: dataB <= 32'b00111011010110000110101100110100;
11'b01100011111: dataB <= 32'b00000101000010010000100010111101;
11'b01100100000: dataB <= 32'b00011101100100110001000110001001;
11'b01100100001: dataB <= 32'b00001001111110011101111010001101;
11'b01100100010: dataB <= 32'b01100110101100001011011000101101;
11'b01100100011: dataB <= 32'b00001101101010011111010001110011;
11'b01100100100: dataB <= 32'b10110000101100011001110101001001;
11'b01100100101: dataB <= 32'b00001000111011111101001001110100;
11'b01100100110: dataB <= 32'b00110110011000100100001100000100;
11'b01100100111: dataB <= 32'b00001001001001001111000101100100;
11'b01100101000: dataB <= 32'b01000111011110111011110101011110;
11'b01100101001: dataB <= 32'b00000111100111101000011010101010;
11'b01100101010: dataB <= 32'b10110101011001000010100010101110;
11'b01100101011: dataB <= 32'b00000101011001011001111010110100;
11'b01100101100: dataB <= 32'b10010101110110101001001001001001;
11'b01100101101: dataB <= 32'b00000011001110011110101101110110;
11'b01100101110: dataB <= 32'b11111010110011011100101111010000;
11'b01100101111: dataB <= 32'b00001010100010100100010010100100;
11'b01100110000: dataB <= 32'b01011100001110011011101000010010;
11'b01100110001: dataB <= 32'b00001000010111111011011010000000;
11'b01100110010: dataB <= 32'b10010101001111101011000100111101;
11'b01100110011: dataB <= 32'b00000100110011011101000100010101;
11'b01100110100: dataB <= 32'b10110000111110100100000101111001;
11'b01100110101: dataB <= 32'b00000101101001010000110111101010;
11'b01100110110: dataB <= 32'b11100101000001110001110110001101;
11'b01100110111: dataB <= 32'b00000000101101110110011011001001;
11'b01100111000: dataB <= 32'b01001110110001111100011110001011;
11'b01100111001: dataB <= 32'b00001001100111011110101110000000;
11'b01100111010: dataB <= 32'b01010111110010011101101011110011;
11'b01100111011: dataB <= 32'b00001110110111100101111011010100;
11'b01100111100: dataB <= 32'b10110110011010001001000111000111;
11'b01100111101: dataB <= 32'b00001001111001101111100001000100;
11'b01100111110: dataB <= 32'b01101110110000100110011101101010;
11'b01100111111: dataB <= 32'b00001101111001111101010001000101;
11'b01101000000: dataB <= 32'b00011011011010010100111111010000;
11'b01101000001: dataB <= 32'b00001011001101001101101111001011;
11'b01101000010: dataB <= 32'b10100000011100011001110000101101;
11'b01101000011: dataB <= 32'b00000101010011001001100101001000;
11'b01101000100: dataB <= 32'b11100001100111001100001010110100;
11'b01101000101: dataB <= 32'b00000111010110100111001111010011;
11'b01101000110: dataB <= 32'b10100110011101011001110000110000;
11'b01101000111: dataB <= 32'b00001101000111001111011010001000;
11'b01101001000: dataB <= 32'b10110010011101111001001010000011;
11'b01101001001: dataB <= 32'b00000111100001101100001010011010;
11'b01101001010: dataB <= 32'b00100001010010110000100001010101;
11'b01101001011: dataB <= 32'b00001010100010110000010010100100;
11'b01101001100: dataB <= 32'b00011000111010010101011011111100;
11'b01101001101: dataB <= 32'b00000111011101111011001010100010;
11'b01101001110: dataB <= 32'b10001100111110000000100010101011;
11'b01101001111: dataB <= 32'b00000111110111010111101110111000;
11'b01101010000: dataB <= 32'b01011000110110001110001011010101;
11'b01101010001: dataB <= 32'b00000010110011100110101100001011;
11'b01101010010: dataB <= 32'b00101100011001100101011000110010;
11'b01101010011: dataB <= 32'b00000111001110100100110000001101;
11'b01101010100: dataB <= 32'b01100000111110100000010110001011;
11'b01101010101: dataB <= 32'b00001011010110101001110001100100;
11'b01101010110: dataB <= 32'b00101010110110101010000100110010;
11'b01101010111: dataB <= 32'b00000101100101001100101110001100;
11'b01101011000: dataB <= 32'b11101111101001001011111001101010;
11'b01101011001: dataB <= 32'b00000000101010001101000010001110;
11'b01101011010: dataB <= 32'b10100000010000100001100100101011;
11'b01101011011: dataB <= 32'b00000100100010011000101001100001;
11'b01101011100: dataB <= 32'b01010110111100101011110101101001;
11'b01101011101: dataB <= 32'b00001010110110101001110110010000;
11'b01101011110: dataB <= 32'b11111100110110011011011011101000;
11'b01101011111: dataB <= 32'b00001111010000111001010011101011;
11'b01101100000: dataB <= 32'b01101100111000001011000011010001;
11'b01101100001: dataB <= 32'b00001110110101110011100010010100;
11'b01101100010: dataB <= 32'b10011100000110111010111110001000;
11'b01101100011: dataB <= 32'b00000101101110010001001101000000;
11'b01101100100: dataB <= 32'b00100011111010110010000101111010;
11'b01101100101: dataB <= 32'b00001010110000101001011010001111;
11'b01101100110: dataB <= 32'b01011110111101010010110111101000;
11'b01101100111: dataB <= 32'b00000111000001000101010001111010;
11'b01101101000: dataB <= 32'b10001101011011011010111100110000;
11'b01101101001: dataB <= 32'b00001011000100101000100100010101;
11'b01101101010: dataB <= 32'b01010101011100011100000001010111;
11'b01101101011: dataB <= 32'b00000110000001011000011101101100;
11'b01101101100: dataB <= 32'b00101101110100110001000110000010;
11'b01101101101: dataB <= 32'b00001100010001110101011111101010;
11'b01101101110: dataB <= 32'b10100000101101000100101001100110;
11'b01101101111: dataB <= 32'b00001100011011110101011110011001;
11'b01101110000: dataB <= 32'b10110001010000001011101000000100;
11'b01101110001: dataB <= 32'b00000011111100101000110011001011;
11'b01101110010: dataB <= 32'b00010011011010100010101001110000;
11'b01101110011: dataB <= 32'b00001101100111111100101110001001;
11'b01101110100: dataB <= 32'b01111101000010100110011101010000;
11'b01101110101: dataB <= 32'b00000010100101001100110011000100;
11'b01101110110: dataB <= 32'b11100101100000010010010101001011;
11'b01101110111: dataB <= 32'b00001100111011101001111010011100;
11'b01101111000: dataB <= 32'b10100010100100001100101000001100;
11'b01101111001: dataB <= 32'b00001100000110100011010001101011;
11'b01101111010: dataB <= 32'b11101010100100001011000011101011;
11'b01101111011: dataB <= 32'b00001010111001111100110101111100;
11'b01101111100: dataB <= 32'b01101100001000101101001001100010;
11'b01101111101: dataB <= 32'b00001000001000010011010001100100;
11'b01101111110: dataB <= 32'b00001101101110110011011000011110;
11'b01101111111: dataB <= 32'b00000110001000100000010110010010;
11'b01110000000: dataB <= 32'b00110111000100110011010010110010;
11'b01110000001: dataB <= 32'b00000111011011100101111010111100;
11'b01110000010: dataB <= 32'b10011111111010001000111000001000;
11'b01110000011: dataB <= 32'b00000011110010011010110010010110;
11'b01110000100: dataB <= 32'b01110110011111011011011110101010;
11'b01110000101: dataB <= 32'b00000111100001011010010010101100;
11'b01110000110: dataB <= 32'b01010100010010011011011000110001;
11'b01110000111: dataB <= 32'b00001001010110111101000001010000;
11'b01110001000: dataB <= 32'b11011001010111011001110111111110;
11'b01110001001: dataB <= 32'b00000101110101011111001000110110;
11'b01110001010: dataB <= 32'b01101110110010100011110111111010;
11'b01110001011: dataB <= 32'b00000100101011010001000011010001;
11'b01110001100: dataB <= 32'b00100100111101011010000110001110;
11'b01110001101: dataB <= 32'b00000000110010101100001010101001;
11'b01110001110: dataB <= 32'b01001111000010000100011100100110;
11'b01110001111: dataB <= 32'b00000111100111011010110001010000;
11'b01110010000: dataB <= 32'b01100001110110101101001100010000;
11'b01110010001: dataB <= 32'b00001111010001101111110011010011;
11'b01110010010: dataB <= 32'b01101100001001100001000101101001;
11'b01110010011: dataB <= 32'b00001011011000110101010001001101;
11'b01110010100: dataB <= 32'b11101010100101000111001100000110;
11'b01110010101: dataB <= 32'b00001111010011111100111001010101;
11'b01110010110: dataB <= 32'b01011111011110011100101110101010;
11'b01110010111: dataB <= 32'b00001010101011010111111011000010;
11'b01110011000: dataB <= 32'b10011000011100001011000000110010;
11'b01110011001: dataB <= 32'b00000110010101010001110000100001;
11'b01110011010: dataB <= 32'b11100111100011001011001011010010;
11'b01110011011: dataB <= 32'b00001000010110101001000111001010;
11'b01110011100: dataB <= 32'b10100000011001000010010001010110;
11'b01110011101: dataB <= 32'b00001011000100010101100101100000;
11'b01110011110: dataB <= 32'b01101010010001011001010111100010;
11'b01110011111: dataB <= 32'b00000100100010100010000110000010;
11'b01110100000: dataB <= 32'b11100101001110000000010010111010;
11'b01110100001: dataB <= 32'b00001000000001100110001010100011;
11'b01110100010: dataB <= 32'b11011000111110100101001101111001;
11'b01110100011: dataB <= 32'b00001001111101111010110110001001;
11'b01110100100: dataB <= 32'b01001101001101011000110010001111;
11'b01110100101: dataB <= 32'b00001001010111100001110010001000;
11'b01110100110: dataB <= 32'b10010110111110100101101011110010;
11'b01110100111: dataB <= 32'b00000011110111100010101000001100;
11'b01110101000: dataB <= 32'b01100100010001111101101001010001;
11'b01110101001: dataB <= 32'b00000110101111100000101100100110;
11'b01110101010: dataB <= 32'b10100000111101110000010101101100;
11'b01110101011: dataB <= 32'b00001100010011110011100101100100;
11'b01110101100: dataB <= 32'b11101000101110010001100101010100;
11'b01110101101: dataB <= 32'b00000011101000001010111110001011;
11'b01110101110: dataB <= 32'b01110101011101001100011000001001;
11'b01110101111: dataB <= 32'b00000000110000001111001110101110;
11'b01110110000: dataB <= 32'b00011000010100001010110100001110;
11'b01110110001: dataB <= 32'b00000010000110010100110001000010;
11'b01110110010: dataB <= 32'b01010111000100110100110100001011;
11'b01110110011: dataB <= 32'b00001011110011110011101001100000;
11'b01110110100: dataB <= 32'b10111000011110010011001001100110;
11'b01110110101: dataB <= 32'b00001111001010111010111111100010;
11'b01110110110: dataB <= 32'b00101000101100001100100011110101;
11'b01110110111: dataB <= 32'b00001111001111111001010010010100;
11'b01110111000: dataB <= 32'b10010000001010101010001100000100;
11'b01110111001: dataB <= 32'b00000101010000010101011000100001;
11'b01110111010: dataB <= 32'b11101111110110010001100111111011;
11'b01110111011: dataB <= 32'b00001010101110101101010010101110;
11'b01110111100: dataB <= 32'b10011110111101001011010110001001;
11'b01110111101: dataB <= 32'b00000100000010001011100101101010;
11'b01110111110: dataB <= 32'b11010011101011000001111100001100;
11'b01110111111: dataB <= 32'b00001000100011100010100000101110;
11'b01111000000: dataB <= 32'b10011101100000100101000011011011;
11'b01111000001: dataB <= 32'b00000011100100010100100101110100;
11'b01111000010: dataB <= 32'b00110101101000010010010011100101;
11'b01111000011: dataB <= 32'b00001100001101111001001011001001;
11'b01111000100: dataB <= 32'b01011100101101001101000111100101;
11'b01111000101: dataB <= 32'b00001101110111111001001001111001;
11'b01111000110: dataB <= 32'b11110011000000001101000110000101;
11'b01111000111: dataB <= 32'b00000110111110100100101111000010;
11'b01111001000: dataB <= 32'b00011001100010010010011001101110;
11'b01111001001: dataB <= 32'b00001011100100110110011001101001;
11'b01111001010: dataB <= 32'b01111010101010111101111100101011;
11'b01111001011: dataB <= 32'b00000001001010001011000011000011;
11'b01111001100: dataB <= 32'b01101011011100001011110100101101;
11'b01111001101: dataB <= 32'b00001110110111110011101110100100;
11'b01111001110: dataB <= 32'b11011110100100011110000111101100;
11'b01111001111: dataB <= 32'b00001010000011100111001101101011;
11'b01111010000: dataB <= 32'b11100100011100001100100011001111;
11'b01111010001: dataB <= 32'b00001100010110111000011110000100;
11'b01111010010: dataB <= 32'b10100000000101000110000110100010;
11'b01111010011: dataB <= 32'b00000110101001010111011101101100;
11'b01111010100: dataB <= 32'b11011001111010101010101011011101;
11'b01111010101: dataB <= 32'b00000100101010010110011001111001;
11'b01111010110: dataB <= 32'b01110110110100110100010011110110;
11'b01111010111: dataB <= 32'b00001001011010101111110010110011;
11'b01111011000: dataB <= 32'b00101011110101100001000110101001;
11'b01111011001: dataB <= 32'b00000100010101011000110110110110;
11'b01111011010: dataB <= 32'b11101110010011001010011101000101;
11'b01111011011: dataB <= 32'b00000101000010010010011010101011;
11'b01111011100: dataB <= 32'b00001100011110001011001000110001;
11'b01111011101: dataB <= 32'b00001010110101111100101000101001;
11'b01111011110: dataB <= 32'b10011101011010111001001010111110;
11'b01111011111: dataB <= 32'b00000110110110100001001001011111;
11'b01111100000: dataB <= 32'b10101010100110011011011001111001;
11'b01111100001: dataB <= 32'b00000100001110010011001110101000;
11'b01111100010: dataB <= 32'b10100100111001000010100101110000;
11'b01111100011: dataB <= 32'b00000001111000100000000110000000;
11'b01111100100: dataB <= 32'b00010001001110000100011010100011;
11'b01111100101: dataB <= 32'b00000110001000011000110100101001;
11'b01111100110: dataB <= 32'b01101011110010110100101011101101;
11'b01111100111: dataB <= 32'b00001111001011110111100011000010;
11'b01111101000: dataB <= 32'b11100000000101000001100100001011;
11'b01111101001: dataB <= 32'b00001100110100110111000001100101;
11'b01111101010: dataB <= 32'b00100100100001110111101010000011;
11'b01111101011: dataB <= 32'b00001111001110111010100001110110;
11'b01111101100: dataB <= 32'b10100101011010011100001101000101;
11'b01111101101: dataB <= 32'b00001001101001100001111010100001;
11'b01111101110: dataB <= 32'b11010100100100001100100001111000;
11'b01111101111: dataB <= 32'b00000111010110011101111000001010;
11'b01111110000: dataB <= 32'b00101101011010111010011011101111;
11'b01111110001: dataB <= 32'b00001001010101101010111110111010;
11'b01111110010: dataB <= 32'b01011000011100110011010010111011;
11'b01111110011: dataB <= 32'b00001000100011011101101000111001;
11'b01111110100: dataB <= 32'b01100000001000111010000101000011;
11'b01111110101: dataB <= 32'b00000010000101010110000101110010;
11'b01111110110: dataB <= 32'b01100111001001010000010101011101;
11'b01111110111: dataB <= 32'b00000101000010011010001010011011;
11'b01111111000: dataB <= 32'b11011001000110101100101111010011;
11'b01111111001: dataB <= 32'b00001100011010110110100001101001;
11'b01111111010: dataB <= 32'b01010001011000110001100010110011;
11'b01111111011: dataB <= 32'b00001010010110101001101101011000;
11'b01111111100: dataB <= 32'b00010111000110111101001100001111;
11'b01111111101: dataB <= 32'b00000101011010011110101000011110;
11'b01111111110: dataB <= 32'b01011100010010001101101001010000;
11'b01111111111: dataB <= 32'b00000110110000011100101101001111;
11'b10000000000: dataB <= 32'b11100000111101000000100101001110;
11'b10000000001: dataB <= 32'b00001100101111111001010101110100;
11'b10000000010: dataB <= 32'b11100100101001110001100110010110;
11'b10000000011: dataB <= 32'b00000010101011001101001110001011;
11'b10000000100: dataB <= 32'b10111001001001011101000111001001;
11'b10000000101: dataB <= 32'b00000001010110010011011011000101;
11'b10000000110: dataB <= 32'b00010000011100001100000100010001;
11'b10000000111: dataB <= 32'b00000000101011010010111000110011;
11'b10000001000: dataB <= 32'b11100011010010011110010101110111;
11'b10000001001: dataB <= 32'b00001001101000110100011000001100;
11'b10000001010: dataB <= 32'b11001110001101100011010011001100;
11'b10000001011: dataB <= 32'b00000101000001011110001001010000;
11'b10000001100: dataB <= 32'b01010110101110010111101010111000;
11'b10000001101: dataB <= 32'b00000111100001101000001110000011;
11'b10000001110: dataB <= 32'b11000101011101000010100010000111;
11'b10000001111: dataB <= 32'b00001000010101101101010100110110;
11'b10000010000: dataB <= 32'b10111010100000110011011101110000;
11'b10000010001: dataB <= 32'b00000111001010101000100111011010;
11'b10000010010: dataB <= 32'b10011111000001101101100100110011;
11'b10000010011: dataB <= 32'b00000001010111110011101001010100;
11'b10000010100: dataB <= 32'b10110101011000111001110110000111;
11'b10000010101: dataB <= 32'b00000001101110010000111011011110;
11'b10000010110: dataB <= 32'b01110001000110100110111101111001;
11'b10000010111: dataB <= 32'b00000010011000010011010110010100;
11'b10000011000: dataB <= 32'b10110100010101001111010010111000;
11'b10000011001: dataB <= 32'b00000110100111100100001100100001;
11'b10000011010: dataB <= 32'b00010111000110100101100010110000;
11'b10000011011: dataB <= 32'b00001011100100100100001100101100;
11'b10000011100: dataB <= 32'b11100000011010100111100010110011;
11'b10000011101: dataB <= 32'b00001111010010010110110101011001;
11'b10000011110: dataB <= 32'b10110001001101001011010111001100;
11'b10000011111: dataB <= 32'b00000010001000001100010000100100;
11'b10000100000: dataB <= 32'b11010100001010111010000101100110;
11'b10000100001: dataB <= 32'b00000101011101100001101001101001;
11'b10000100010: dataB <= 32'b11101110101001111111100110110110;
11'b10000100011: dataB <= 32'b00001011100010110110011010001010;
11'b10000100100: dataB <= 32'b10010011000011000111000110010000;
11'b10000100101: dataB <= 32'b00000001101011100110110001111100;
11'b10000100110: dataB <= 32'b11001110110110010111100111111001;
11'b10000100111: dataB <= 32'b00001011000111001110001110011011;
11'b10000101000: dataB <= 32'b10000010111111000101110001010010;
11'b10000101001: dataB <= 32'b00000100110010101111010010010100;
11'b10000101010: dataB <= 32'b00111101001101010010101110101001;
11'b10000101011: dataB <= 32'b00000101010110001101010000111100;
11'b10000101100: dataB <= 32'b01011010010010001110011011011000;
11'b10000101101: dataB <= 32'b00001101001101111000100001101010;
11'b10000101110: dataB <= 32'b01111010101000100100110100110010;
11'b10000101111: dataB <= 32'b00001010110111011011001111000010;
11'b10000110000: dataB <= 32'b10001000100001001001100010100101;
11'b10000110001: dataB <= 32'b00000001010101001101011001111010;
11'b10000110010: dataB <= 32'b10001111100101100011101000101110;
11'b10000110011: dataB <= 32'b00001010101010010100000100100110;
11'b10000110100: dataB <= 32'b00101101000100100010001111001010;
11'b10000110101: dataB <= 32'b00001011010010100100111111110101;
11'b10000110110: dataB <= 32'b10010010101001101011001100101100;
11'b10000110111: dataB <= 32'b00000111010111100111011000010010;
11'b10000111000: dataB <= 32'b11011100110101010101111000010100;
11'b10000111001: dataB <= 32'b00001100011100000010111100010011;
11'b10000111010: dataB <= 32'b10100111011110001011110001101010;
11'b10000111011: dataB <= 32'b00000100010011011011001100100110;
11'b10000111100: dataB <= 32'b11111000101010010010010110101000;
11'b10000111101: dataB <= 32'b00000101100001110000010001001001;
11'b10000111110: dataB <= 32'b11000010111100110101110101110111;
11'b10000111111: dataB <= 32'b00001010000110100000010010111100;
11'b10001000000: dataB <= 32'b01010000110111110100010001101011;
11'b10001000001: dataB <= 32'b00000111000001010000001011000100;
11'b10001000010: dataB <= 32'b11101100110110000011000010100101;
11'b10001000011: dataB <= 32'b00000100101100111100111100110010;
11'b10001000100: dataB <= 32'b10010011010110010111101100011100;
11'b10001000101: dataB <= 32'b00001011010001111101000101011111;
11'b10001000110: dataB <= 32'b00101100100101001010000111101000;
11'b10001000111: dataB <= 32'b00001010101101011110101001000010;
11'b10001001000: dataB <= 32'b00001111001101101110011101111010;
11'b10001001001: dataB <= 32'b00000001101110110101000100101110;
11'b10001001010: dataB <= 32'b01000100111101000110000001110101;
11'b10001001011: dataB <= 32'b00000010111011000011010001001100;
11'b10001001100: dataB <= 32'b00100100110000001101011110110101;
11'b10001001101: dataB <= 32'b00000001010101000101001001101011;
11'b10001001110: dataB <= 32'b10100011001110010010101001100001;
11'b10001001111: dataB <= 32'b00001101000111010000010000111100;
11'b10001010000: dataB <= 32'b00101101011100110110011001111010;
11'b10001010001: dataB <= 32'b00001011001011110110101100001101;
11'b10001010010: dataB <= 32'b00100011010010100010000111100111;
11'b10001010011: dataB <= 32'b00001101010101010101000011000111;
11'b10001010100: dataB <= 32'b10001001000110110011101000001101;
11'b10001010101: dataB <= 32'b00001000010010010111000111101101;
11'b10001010110: dataB <= 32'b01011110111100010101110111010101;
11'b10001010111: dataB <= 32'b00000111100110101010001110011100;
11'b10001011000: dataB <= 32'b10010100110100110100011011010011;
11'b10001011001: dataB <= 32'b00000101111010100111100101111011;
11'b10001011010: dataB <= 32'b11100100001110100101000100110001;
11'b10001011011: dataB <= 32'b00001011011101101101011010110001;
11'b10001011100: dataB <= 32'b01001111011110000111101000110111;
11'b10001011101: dataB <= 32'b00000101111110011101011001100110;
11'b10001011110: dataB <= 32'b01011111010001111110100100110100;
11'b10001011111: dataB <= 32'b00001011001010111010101100001011;
11'b10001100000: dataB <= 32'b10011010000101101011000100001000;
11'b10001100001: dataB <= 32'b00001000000001101000001101111000;
11'b10001100010: dataB <= 32'b01011100100101100111101000111001;
11'b10001100011: dataB <= 32'b00001010100010110000011010001011;
11'b10001100100: dataB <= 32'b11000011000101011010000100000011;
11'b10001100101: dataB <= 32'b00000111010100100111011100010101;
11'b10001100110: dataB <= 32'b10111100111001000010011101010100;
11'b10001100111: dataB <= 32'b00001000001010101100101111100011;
11'b10001101000: dataB <= 32'b00011111000001011101010100010000;
11'b10001101001: dataB <= 32'b00000000110001101001110101001100;
11'b10001101010: dataB <= 32'b01101101100101011001001000000110;
11'b10001101011: dataB <= 32'b00000010001001010010101110110111;
11'b10001101100: dataB <= 32'b10101111010110000111001011111101;
11'b10001101101: dataB <= 32'b00000000110011001111001110001100;
11'b10001101110: dataB <= 32'b10111010100100100110010001010011;
11'b10001101111: dataB <= 32'b00001000100111101110010101000000;
11'b10001110000: dataB <= 32'b00010110111110010101110011001100;
11'b10001110001: dataB <= 32'b00001101100111101110010100110011;
11'b10001110010: dataB <= 32'b10101000011101110111100010001111;
11'b10001110011: dataB <= 32'b00001110011000011000101101110001;
11'b10001110100: dataB <= 32'b10101101011001010010111000001100;
11'b10001110101: dataB <= 32'b00000011100100010110000100100011;
11'b10001110110: dataB <= 32'b11100000000111001010111000000101;
11'b10001110111: dataB <= 32'b00000010111010011001100110001001;
11'b10001111000: dataB <= 32'b00110000110101001111010101110101;
11'b10001111001: dataB <= 32'b00001101100110111100101110011011;
11'b10001111010: dataB <= 32'b10010010111010010111100110001111;
11'b10001111011: dataB <= 32'b00000011000111101000111001110100;
11'b10001111100: dataB <= 32'b00010010101001100111100101111000;
11'b10001111101: dataB <= 32'b00001100101010011010000110011100;
11'b10001111110: dataB <= 32'b11000100100110100110100001001100;
11'b10001111111: dataB <= 32'b00000100001111101001011010001100;
11'b10010000000: dataB <= 32'b01110111100101101010011111001111;
11'b10010000001: dataB <= 32'b00000100010011001010111101000011;
11'b10010000010: dataB <= 32'b00100010010001101110011001011010;
11'b10010000011: dataB <= 32'b00001101110001111100110110000010;
11'b10010000100: dataB <= 32'b01111101000000011011100100001111;
11'b10010000101: dataB <= 32'b00001001011000011001001011010011;
11'b10010000110: dataB <= 32'b10001110010001101001000101000010;
11'b10010000111: dataB <= 32'b00000000110000001001001010001010;
11'b10010001000: dataB <= 32'b01001001010101101011001000101110;
11'b10010001001: dataB <= 32'b00001011001101100000000100001101;
11'b10010001010: dataB <= 32'b01101011001100111001001111010000;
11'b10010001011: dataB <= 32'b00001010110100100101000011011110;
11'b10010001100: dataB <= 32'b01011000100001111010111101010000;
11'b10010001101: dataB <= 32'b00000101110110100001011100101001;
11'b10010001110: dataB <= 32'b10011110110101000101000111010011;
11'b10010001111: dataB <= 32'b00001001011110000100100100100010;
11'b10010010000: dataB <= 32'b01100001100010001011110011000110;
11'b10010010001: dataB <= 32'b00000011110000011001001000001101;
11'b10010010010: dataB <= 32'b01111010111110100010101000000111;
11'b10010010011: dataB <= 32'b00001000100001111000100001101001;
11'b10010010100: dataB <= 32'b10000100100100100100110100110100;
11'b10010010101: dataB <= 32'b00001100001001101000010110101101;
11'b10010010110: dataB <= 32'b01010010101011100101110011000111;
11'b10010010111: dataB <= 32'b00001001100001011100000110111101;
11'b10010011000: dataB <= 32'b11101111000010010011000101000010;
11'b10010011001: dataB <= 32'b00000101101010111101010001001001;
11'b10010011010: dataB <= 32'b11001111001101100111101001011110;
11'b10010011011: dataB <= 32'b00001010110011111001011100110110;
11'b10010011100: dataB <= 32'b10110000110001100001101001001001;
11'b10010011101: dataB <= 32'b00001011001111100010101101011001;
11'b10010011110: dataB <= 32'b11001100111101001101111011011101;
11'b10010011111: dataB <= 32'b00000010001001110011010100010100;
11'b10010100000: dataB <= 32'b11001000101000101101000001010000;
11'b10010100001: dataB <= 32'b00000001010110000010111001001011;
11'b10010100010: dataB <= 32'b11100110110100001011111101011010;
11'b10010100011: dataB <= 32'b00000000101111000100110001111010;
11'b10010100100: dataB <= 32'b10011111001110100010111100100100;
11'b10010100101: dataB <= 32'b00001110101100011010001000111011;
11'b10010100110: dataB <= 32'b10100111100100011101000111111011;
11'b10010100111: dataB <= 32'b00001011101101111000111100001011;
11'b10010101000: dataB <= 32'b10011111010010110010111001001000;
11'b10010101001: dataB <= 32'b00001011111000010100111010010111;
11'b10010101010: dataB <= 32'b11001000110110110100001000101101;
11'b10010101011: dataB <= 32'b00000111110010010110111111001110;
11'b10010101100: dataB <= 32'b11011110111100001100010110010100;
11'b10010101101: dataB <= 32'b00001001100111110010011010010100;
11'b10010101110: dataB <= 32'b10010110101100110011011010010101;
11'b10010101111: dataB <= 32'b00000100011000011111101001111011;
11'b10010110000: dataB <= 32'b10101110010110001101100100101111;
11'b10010110001: dataB <= 32'b00001000011110100111100011001010;
11'b10010110010: dataB <= 32'b11001011001101011111100111010111;
11'b10010110011: dataB <= 32'b00000011011011011001010101000101;
11'b10010110100: dataB <= 32'b00011011001101011110010011110001;
11'b10010110101: dataB <= 32'b00001011101101111101000100011010;
11'b10010110110: dataB <= 32'b11100100000101111010110110000110;
11'b10010110111: dataB <= 32'b00001011000010110010011010100000;
11'b10010111000: dataB <= 32'b10100000100100111111000111011001;
11'b10010111001: dataB <= 32'b00001101000101110110101010010011;
11'b10010111010: dataB <= 32'b01000010101101110001110110100001;
11'b10010111011: dataB <= 32'b00000110010011100001100000001100;
11'b10010111100: dataB <= 32'b11111101001101011001111011111000;
11'b10010111101: dataB <= 32'b00001001001010101110111011100100;
11'b10010111110: dataB <= 32'b10011111000001001100110100001101;
11'b10010111111: dataB <= 32'b00000000101011011101111001001011;
11'b10011000000: dataB <= 32'b10100101101110000000111001100111;
11'b10011000001: dataB <= 32'b00000011100101010110100110000111;
11'b10011000010: dataB <= 32'b11101011011101011110111000111110;
11'b10011000011: dataB <= 32'b00000000101101001110111110000100;
11'b10011000100: dataB <= 32'b01111100111100001101000001001110;
11'b10011000101: dataB <= 32'b00001010001000110100100001110000;
11'b10011000110: dataB <= 32'b01011000110101111101110011101001;
11'b10011000111: dataB <= 32'b00001110101100110100100000111010;
11'b10011001000: dataB <= 32'b11101100101001000111010010101011;
11'b10011001001: dataB <= 32'b00001100011100011100101010010001;
11'b10011001010: dataB <= 32'b01100111100001100010011000101100;
11'b10011001011: dataB <= 32'b00000110000010100010000100101010;
11'b10011001100: dataB <= 32'b00101010001011010011111010000110;
11'b10011001101: dataB <= 32'b00000001010101010001011110100010;
11'b10011001110: dataB <= 32'b10110011000100100110010100110011;
11'b10011001111: dataB <= 32'b00001111001100111101000110100011;
11'b10011010000: dataB <= 32'b01010110110001101111100110101110;
11'b10011010001: dataB <= 32'b00000101000100101001000001101100;
11'b10011010010: dataB <= 32'b01010110011100111111000100110101;
11'b10011010011: dataB <= 32'b00001101101110100100000110010100;
11'b10011010100: dataB <= 32'b11001100010010000110110010000111;
11'b10011010101: dataB <= 32'b00000100101101100011100010000100;
11'b10011010110: dataB <= 32'b10101111110001111010001111010101;
11'b10011010111: dataB <= 32'b00000011110000001100101101001010;
11'b10011011000: dataB <= 32'b01101100010101010101110111011010;
11'b10011011001: dataB <= 32'b00001100110101111101001110010010;
11'b10011011010: dataB <= 32'b01111011010100100010100100101101;
11'b10011011011: dataB <= 32'b00000111011001010111000011010100;
11'b10011011100: dataB <= 32'b11011000001010010001001000000001;
11'b10011011101: dataB <= 32'b00000001001010001000110110011010;
11'b10011011110: dataB <= 32'b11000111000101110011001001001111;
11'b10011011111: dataB <= 32'b00001011101111101100001000001011;
11'b10011100000: dataB <= 32'b01100111010101100000101110110110;
11'b10011100001: dataB <= 32'b00001001110110100011000110110111;
11'b10011100010: dataB <= 32'b10011110011110000010111100110100;
11'b10011100011: dataB <= 32'b00000100110100011011011101010000;
11'b10011100100: dataB <= 32'b10100000110100111100010110110011;
11'b10011100101: dataB <= 32'b00000110111110001100010000111001;
11'b10011100110: dataB <= 32'b11011001100010001100000101100011;
11'b10011100111: dataB <= 32'b00000011101100010111000000001011;
11'b10011101000: dataB <= 32'b01111001010010110011001001101000;
11'b10011101001: dataB <= 32'b00001011100010111100110110001001;
11'b10011101010: dataB <= 32'b11001100010000100011100011110001;
11'b10011101011: dataB <= 32'b00001100101100110000100010010101;
11'b10011101100: dataB <= 32'b11011000100011001110110101000100;
11'b10011101101: dataB <= 32'b00001100100100101000000110101101;
11'b10011101110: dataB <= 32'b10101101001010011011011000000001;
11'b10011101111: dataB <= 32'b00000110101001110111100101100001;
11'b10011110000: dataB <= 32'b10001110111100111111000110111110;
11'b10011110001: dataB <= 32'b00001001110101110011101100010101;
11'b10011110010: dataB <= 32'b01110010111110000001101010001010;
11'b10011110011: dataB <= 32'b00001011010001100110110001111001;
11'b10011110100: dataB <= 32'b10001110110000111101001000011110;
11'b10011110101: dataB <= 32'b00000011100101101101100000010011;
11'b10011110110: dataB <= 32'b00001110011000100100000001101011;
11'b10011110111: dataB <= 32'b00000000110000000100100101010011;
11'b10011111000: dataB <= 32'b11101000111100010010011010111101;
11'b10011111001: dataB <= 32'b00000001001010001000011110000010;
11'b10011111010: dataB <= 32'b11011101001110101011011110001000;
11'b10011111011: dataB <= 32'b00001110110001100100001001000010;
11'b10011111100: dataB <= 32'b00011111100100010011110101111010;
11'b10011111101: dataB <= 32'b00001011110000110111010000010010;
11'b10011111110: dataB <= 32'b10011011001111000011101010101001;
11'b10011111111: dataB <= 32'b00001001111010010110110001101111;
11'b10100000000: dataB <= 32'b10001100100110101100111001001110;
11'b10100000001: dataB <= 32'b00000111010001011000110110100111;
11'b10100000010: dataB <= 32'b11011110111100001010110101110011;
11'b10100000011: dataB <= 32'b00001011001001111000101110001100;
11'b10100000100: dataB <= 32'b10011010101001000010101001010110;
11'b10100000101: dataB <= 32'b00000010110100010111100110000011;
11'b10100000110: dataB <= 32'b10110100100001111101100101001100;
11'b10100000111: dataB <= 32'b00000101011110100001100111011011;
11'b10100001000: dataB <= 32'b11001000111100110110110101110110;
11'b10100001001: dataB <= 32'b00000001010110010101001100110100;
11'b10100001010: dataB <= 32'b11011001001001000101100011101110;
11'b10100001011: dataB <= 32'b00001100010000111001011000111000;
11'b10100001100: dataB <= 32'b10110000001110001010111000000101;
11'b10100001101: dataB <= 32'b00001101100101111000101011001001;
11'b10100001110: dataB <= 32'b11100100101000011110000101011000;
11'b10100001111: dataB <= 32'b00001110101010111010111110010011;
11'b10100010000: dataB <= 32'b11001000011010010001111001100010;
11'b10100010001: dataB <= 32'b00000101110001011011011100001010;
11'b10100010010: dataB <= 32'b00110111100101111001011010011010;
11'b10100010011: dataB <= 32'b00001010001100101111000111001110;
11'b10100010100: dataB <= 32'b11011111000001000100000100101011;
11'b10100010101: dataB <= 32'b00000010000110010011110001011010;
11'b10100010110: dataB <= 32'b10011101101110100001001011001001;
11'b10100010111: dataB <= 32'b00000110000011011100100001010111;
11'b10100011000: dataB <= 32'b11100011100000111110000101111110;
11'b10100011001: dataB <= 32'b00000001101000010000110001111100;
11'b10100011010: dataB <= 32'b01111101010100001011110010001001;
11'b10100011011: dataB <= 32'b00001011101010111000110110100000;
11'b10100011100: dataB <= 32'b10011010110001100101100101100110;
11'b10100011101: dataB <= 32'b00001110110010111000110101011001;
11'b10100011110: dataB <= 32'b00110000110100100110010100000111;
11'b10100011111: dataB <= 32'b00001001011110100000101010101010;
11'b10100100000: dataB <= 32'b10011111100101111010001001001101;
11'b10100100001: dataB <= 32'b00001001000010101110001001000001;
11'b10100100010: dataB <= 32'b10110100010111001101001011101000;
11'b10100100011: dataB <= 32'b00000000101111001101001110111010;
11'b10100100100: dataB <= 32'b00110001010000001101000100010000;
11'b10100100101: dataB <= 32'b00001111010001111011011110101100;
11'b10100100110: dataB <= 32'b00011000101000111111000111001101;
11'b10100100111: dataB <= 32'b00000111100010101001001001101100;
11'b10100101000: dataB <= 32'b10011110011000011110000011110010;
11'b10100101001: dataB <= 32'b00001101010010110000001110001100;
11'b10100101010: dataB <= 32'b11010110000101100110100100000100;
11'b10100101011: dataB <= 32'b00000101001010011101100001110100;
11'b10100101100: dataB <= 32'b00100011111010010010011101111010;
11'b10100101101: dataB <= 32'b00000100001101010000100001100010;
11'b10100101110: dataB <= 32'b10110010100000111101000101011001;
11'b10100101111: dataB <= 32'b00001011011000110111100010101010;
11'b10100110000: dataB <= 32'b01110101101000111001100101001010;
11'b10100110001: dataB <= 32'b00000101111000010110111011001101;
11'b10100110010: dataB <= 32'b01100100001010110001101010100010;
11'b10100110011: dataB <= 32'b00000010100101001100100110100011;
11'b10100110100: dataB <= 32'b01001000110010000010111001010000;
11'b10100110101: dataB <= 32'b00001011010010110110010100010010;
11'b10100110110: dataB <= 32'b10100011011010010000101101011011;
11'b10100110111: dataB <= 32'b00001000010111100011000110000111;
11'b10100111000: dataB <= 32'b01100100100010010011001011010111;
11'b10100111001: dataB <= 32'b00000100010001010111011010000000;
11'b10100111010: dataB <= 32'b11100010110100111011010110010001;
11'b10100111011: dataB <= 32'b00000011111100010110000101011000;
11'b10100111100: dataB <= 32'b01010101011010001100001000000010;
11'b10100111101: dataB <= 32'b00000100101010010110111000010010;
11'b10100111110: dataB <= 32'b10110011100110111011111011001010;
11'b10100111111: dataB <= 32'b00001101100110111011001110101001;
11'b10101000000: dataB <= 32'b00010110000100101010010011101110;
11'b10101000001: dataB <= 32'b00001101010000110100101101111110;
11'b10101000010: dataB <= 32'b00011110011110011111100111100010;
11'b10101000011: dataB <= 32'b00001110101000110010010010001110;
11'b10101000100: dataB <= 32'b01101011010110011011111010100010;
11'b10101000101: dataB <= 32'b00001000001000101101110110000001;
11'b10101000110: dataB <= 32'b00010000110000011110000011111100;
11'b10101000111: dataB <= 32'b00001000110110100111111000001100;
11'b10101001000: dataB <= 32'b10110001001110100001101011001100;
11'b10101001001: dataB <= 32'b00001010010100101000111010100001;
11'b10101001010: dataB <= 32'b01010010100100101100000101011110;
11'b10101001011: dataB <= 32'b00000110000011100111101000100010;
11'b10101001100: dataB <= 32'b10010110001100101011000011000110;
11'b10101001101: dataB <= 32'b00000000101010001100010001011010;
11'b10101001110: dataB <= 32'b00101001000100101001010111111110;
11'b10101001111: dataB <= 32'b00000010100101010000010010010011;
11'b10101010000: dataB <= 32'b00011011001010110011111111001110;
11'b10101010001: dataB <= 32'b00001101110110101110010001010010;
11'b10101010010: dataB <= 32'b00010111100100011010100011110111;
11'b10101010011: dataB <= 32'b00001011010011110001100000110001;
11'b10101010100: dataB <= 32'b00011001001011000100011011101100;
11'b10101010101: dataB <= 32'b00000111111011011010101100111111;
11'b10101010110: dataB <= 32'b10010010010110100101011001001111;
11'b10101010111: dataB <= 32'b00000111010001011010110001111111;
11'b10101011000: dataB <= 32'b00011110111100100001100101010001;
11'b10101011001: dataB <= 32'b00001100001100111011000001111101;
11'b10101011010: dataB <= 32'b10011110100101011001110111110111;
11'b10101011011: dataB <= 32'b00000010010000010001011010000011;
11'b10101011100: dataB <= 32'b10111000110101101101010101101010;
11'b10101011101: dataB <= 32'b00000010111011011001100011010100;
11'b10101011110: dataB <= 32'b11001010101000010101100100110100;
11'b10101011111: dataB <= 32'b00000000110000010011000100101011;
endcase
end
assign doA = dataA;
assign doB = dataB;
endmodule
