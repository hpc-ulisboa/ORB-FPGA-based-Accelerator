module rams_sp_rom1_8_sec (clk, enA, enB, addrA, addrB, doA, doB);
input clk;
input enA, enB;
input [11:0] addrA, addrB;
output [31:0] doA, doB;
(*rom_style = "block" *) reg [2751:0] dataA, dataB;
always @(posedge clk)
begin
if (enA)
case(addrA)
12'b000000000000: dataA <= 32'b00000111001100111111000001110111;
12'b000000000001: dataA <= 32'b00001011010000010011000111110100;
12'b000000000010: dataA <= 32'b00001100010011010110101010011001;
12'b000000000011: dataA <= 32'b00001110000111101010010000110010;
12'b000000000100: dataA <= 32'b10010111111010100010000111100111;
12'b000000000101: dataA <= 32'b00001111001100101010110010000111;
12'b000000000110: dataA <= 32'b00010011001101101110100110110101;
12'b000000000111: dataA <= 32'b00000110101010010000100011110101;
12'b000000001000: dataA <= 32'b00000100100010110011001000101011;
12'b000000001001: dataA <= 32'b00000100110110000101011011010010;
12'b000000001010: dataA <= 32'b11011111001011110100101011110011;
12'b000000001011: dataA <= 32'b00001011001101000010110110100100;
12'b000000001100: dataA <= 32'b01011010110110001001110110000011;
12'b000000001101: dataA <= 32'b00000011001100110000100110010011;
12'b000000001110: dataA <= 32'b10101111100101110001010100000011;
12'b000000001111: dataA <= 32'b00001110101001011000101010010111;
12'b000000010000: dataA <= 32'b10101111010011000101101001110010;
12'b000000010001: dataA <= 32'b00000000110010101100111001010110;
12'b000000010010: dataA <= 32'b00100010001011001001000011100011;
12'b000000010011: dataA <= 32'b00001011001011111000100010110001;
12'b000000010100: dataA <= 32'b01001101001110100010001001100001;
12'b000000010101: dataA <= 32'b00001010001011010000100100100110;
12'b000000010110: dataA <= 32'b00011011010101111100001010101110;
12'b000000010111: dataA <= 32'b00001111001010000100110110010101;
12'b000000011000: dataA <= 32'b01000100101011011110011111010100;
12'b000000011001: dataA <= 32'b00001001101100110000101110100010;
12'b000000011010: dataA <= 32'b10010001011101001011101011001100;
12'b000000011011: dataA <= 32'b00000001101000001110001101011111;
12'b000000011100: dataA <= 32'b00100011011011001100000001010000;
12'b000000011101: dataA <= 32'b00001111010001011111000101010110;
12'b000000011110: dataA <= 32'b00011001111011101101111011110110;
12'b000000011111: dataA <= 32'b00001101110101100111010111000111;
12'b000000100000: dataA <= 32'b01000111100000111111001011010001;
12'b000000100001: dataA <= 32'b00001100001000100110011110011110;
12'b000000100010: dataA <= 32'b10100111010101110100111001110001;
12'b000000100011: dataA <= 32'b00000100011000011011001110001110;
12'b000000100100: dataA <= 32'b11100110010111110010110011101011;
12'b000000100101: dataA <= 32'b00000101111110011111100001111001;
12'b000000100110: dataA <= 32'b10001110101111110011000111101110;
12'b000000100111: dataA <= 32'b00001110110111010101011110001010;
12'b000000101000: dataA <= 32'b01010001000101111001110010001000;
12'b000000101001: dataA <= 32'b00001000111000011001011101110100;
12'b000000101010: dataA <= 32'b01101011010011110101001011110010;
12'b000000101011: dataA <= 32'b00001100010001011001000011000110;
12'b000000101100: dataA <= 32'b10101011001000111101111101110011;
12'b000000101101: dataA <= 32'b00001100000111010100001101000101;
12'b000000101110: dataA <= 32'b11101000001011101010011010101000;
12'b000000101111: dataA <= 32'b00001101010010001101000101101010;
12'b000000110000: dataA <= 32'b00100011001101010100000001001111;
12'b000000110001: dataA <= 32'b00000101001101001010101110011110;
12'b000000110010: dataA <= 32'b11100011011001010001111011100010;
12'b000000110011: dataA <= 32'b00001011010110010001011110110101;
12'b000000110100: dataA <= 32'b10011001101011001100101010010001;
12'b000000110101: dataA <= 32'b00001011001001010100101010100111;
12'b000000110110: dataA <= 32'b10011100010100110010010010100101;
12'b000000110111: dataA <= 32'b00001100111010011011010101010001;
12'b000000111000: dataA <= 32'b11110000110011001001000110100110;
12'b000000111001: dataA <= 32'b00001001010010011011001000010011;
12'b000000111010: dataA <= 32'b00011011011011000010110010001011;
12'b000000111011: dataA <= 32'b00001010001010110000001111011101;
12'b000000111100: dataA <= 32'b01100000100001101011010011101100;
12'b000000111101: dataA <= 32'b00000001001001000110011110110010;
12'b000000111110: dataA <= 32'b10101011000011001001111010100010;
12'b000000111111: dataA <= 32'b00000010111010100001000000011101;
12'b000001000000: dataA <= 32'b11001010111110001010010110000111;
12'b000001000001: dataA <= 32'b00000010101001011110001011110011;
12'b000001000010: dataA <= 32'b01001110011001000010110010100111;
12'b000001000011: dataA <= 32'b00001010110111010101010000010010;
12'b000001000100: dataA <= 32'b11110000011001111101010001110101;
12'b000001000101: dataA <= 32'b00000011110011100100111110010010;
12'b000001000110: dataA <= 32'b10000100101011011110010010011001;
12'b000001000111: dataA <= 32'b00001011110010100101000101010010;
12'b000001001000: dataA <= 32'b10000101000011000011000011001101;
12'b000001001001: dataA <= 32'b00001001101100010000110110100011;
12'b000001001010: dataA <= 32'b00011111001100101110100011110110;
12'b000001001011: dataA <= 32'b00001010111110100001101111110101;
12'b000001001100: dataA <= 32'b00101010001010000001110100100110;
12'b000001001101: dataA <= 32'b00000001100111110100010101111001;
12'b000001001110: dataA <= 32'b00010000001101100010101011100110;
12'b000001001111: dataA <= 32'b00001101010110001111010101101010;
12'b000001010000: dataA <= 32'b10100001001001010111010111011011;
12'b000001010001: dataA <= 32'b00001100101111100110111010101100;
12'b000001010010: dataA <= 32'b00011001011101010110011100110111;
12'b000001010011: dataA <= 32'b00001011100101100110010100011110;
12'b000001010100: dataA <= 32'b00000000000000101100010100101111;
12'b000001010101: dataA <= 32'b00000000000000000000000000000000;
12'b000001010110: dataA <= 32'b01001001010101001111010010011010;
12'b000001010111: dataA <= 32'b00001011001111010011001011110011;
12'b000001011000: dataA <= 32'b10001000011011011101111011011000;
12'b000001011001: dataA <= 32'b00001101000100100110001100101010;
12'b000001011010: dataA <= 32'b10011101111010010001110110100111;
12'b000001011011: dataA <= 32'b00001110101001101000101110011111;
12'b000001011100: dataA <= 32'b01010101010010000110100111010101;
12'b000001011101: dataA <= 32'b00000110001010001100101011110100;
12'b000001011110: dataA <= 32'b11000010101110101010111000001011;
12'b000001011111: dataA <= 32'b00000101110111000111100011000001;
12'b000001100000: dataA <= 32'b10011111001011110011111011110001;
12'b000001100001: dataA <= 32'b00001011001100000011000010100100;
12'b000001100010: dataA <= 32'b01011010110101111001110101000100;
12'b000001100011: dataA <= 32'b00000011001110101100011110010011;
12'b000001100100: dataA <= 32'b10110011011101100001010011000101;
12'b000001100101: dataA <= 32'b00001101100110010110101110101111;
12'b000001100110: dataA <= 32'b11110001001011001101001001110001;
12'b000001100111: dataA <= 32'b00000000110101101100110101100110;
12'b000001101000: dataA <= 32'b11011110001010111000100010100101;
12'b000001101001: dataA <= 32'b00001010101010110110010110100000;
12'b000001101010: dataA <= 32'b11001111010110010001111000000001;
12'b000001101011: dataA <= 32'b00001001101010001110101100110110;
12'b000001101100: dataA <= 32'b00011101010101111100001010101101;
12'b000001101101: dataA <= 32'b00001110001000000100111110011101;
12'b000001101110: dataA <= 32'b00000010110111101101111111010010;
12'b000001101111: dataA <= 32'b00001001001011101110100110011010;
12'b000001110000: dataA <= 32'b10010101100101001011111010101011;
12'b000001110001: dataA <= 32'b00000000101011001010010101101111;
12'b000001110010: dataA <= 32'b01100101011011000011100001110010;
12'b000001110011: dataA <= 32'b00001111001110011111000101100110;
12'b000001110100: dataA <= 32'b10011111111011110101001100010100;
12'b000001110101: dataA <= 32'b00001110010011101001010011011110;
12'b000001110110: dataA <= 32'b00001011101101001111011011010000;
12'b000001110111: dataA <= 32'b00001011000110100010011110101110;
12'b000001111000: dataA <= 32'b10101001010001110100111001110001;
12'b000001111001: dataA <= 32'b00000101011001011101001110011110;
12'b000001111010: dataA <= 32'b11100010010011101010000011001101;
12'b000001111011: dataA <= 32'b00000111011110100011011101101001;
12'b000001111100: dataA <= 32'b10001100110111101010010111101110;
12'b000001111101: dataA <= 32'b00001111010100011001100010000010;
12'b000001111110: dataA <= 32'b01010001001101101001110001001010;
12'b000001111111: dataA <= 32'b00001001111000011101011101110100;
12'b000010000000: dataA <= 32'b11101101001111110100101011110000;
12'b000010000001: dataA <= 32'b00001100001111011001000111010101;
12'b000010000010: dataA <= 32'b00101011000101001110011101110001;
12'b000010000011: dataA <= 32'b00001011000101010000010001010110;
12'b000010000100: dataA <= 32'b11100010000111011001101001100111;
12'b000010000101: dataA <= 32'b00001101001111001101001101100010;
12'b000010000110: dataA <= 32'b11100101001101010100010001010001;
12'b000010000111: dataA <= 32'b00000101001110001000110110101101;
12'b000010001000: dataA <= 32'b01100101011001000010001010000001;
12'b000010001001: dataA <= 32'b00001011110100010101100111000101;
12'b000010001010: dataA <= 32'b01011101101111001100001010010000;
12'b000010001011: dataA <= 32'b00001010001000010010101110111111;
12'b000010001100: dataA <= 32'b11011000010100101010110001101000;
12'b000010001101: dataA <= 32'b00001101011000011101010101000001;
12'b000010001110: dataA <= 32'b01101110101010111000110101100111;
12'b000010001111: dataA <= 32'b00001001010010011011001000010100;
12'b000010010000: dataA <= 32'b10011101011010111010010001101101;
12'b000010010001: dataA <= 32'b00001001101001101010001011100100;
12'b000010010010: dataA <= 32'b00011100100101101011010011101110;
12'b000010010011: dataA <= 32'b00000000101100000100100110100010;
12'b000010010100: dataA <= 32'b00101010111110111001011001000001;
12'b000010010101: dataA <= 32'b00000011111100100001000000101110;
12'b000010010110: dataA <= 32'b00001101000110000010010101001000;
12'b000010010111: dataA <= 32'b00000010001011011010001111110011;
12'b000010011000: dataA <= 32'b00001010100000111011010001101001;
12'b000010011001: dataA <= 32'b00001011110110010111010100001011;
12'b000010011010: dataA <= 32'b11101010010010000101010010010111;
12'b000010011011: dataA <= 32'b00000100010101100100111110001010;
12'b000010011100: dataA <= 32'b11000010110111101101110011011011;
12'b000010011101: dataA <= 32'b00001011110000100101000101001010;
12'b000010011110: dataA <= 32'b01000111001010111010100011001111;
12'b000010011111: dataA <= 32'b00001001001011010000111110100011;
12'b000010100000: dataA <= 32'b10011111001100111111000100111000;
12'b000010100001: dataA <= 32'b00001011111100100101101011110100;
12'b000010100010: dataA <= 32'b01100100000101110010000011101000;
12'b000010100011: dataA <= 32'b00000001001010101110001101101001;
12'b000010100100: dataA <= 32'b00001100010101011010111010100101;
12'b000010100101: dataA <= 32'b00001101110100010001011101011010;
12'b000010100110: dataA <= 32'b01100001001001101111101000011011;
12'b000010100111: dataA <= 32'b00001100101101100110110110101100;
12'b000010101000: dataA <= 32'b10011101011101100110101101010101;
12'b000010101001: dataA <= 32'b00001010100011100000010100101110;
12'b000010101010: dataA <= 32'b00000000000000101100110100110000;
12'b000010101011: dataA <= 32'b00000000000000000000000000000000;
12'b000010101100: dataA <= 32'b10001011011101100111100011111100;
12'b000010101101: dataA <= 32'b00001010101110010101010011110010;
12'b000010101110: dataA <= 32'b01000110100011101101011100010110;
12'b000010101111: dataA <= 32'b00001011100011100000001000100011;
12'b000010110000: dataA <= 32'b01100011111010001001110101101000;
12'b000010110001: dataA <= 32'b00001110000111100110101010110111;
12'b000010110010: dataA <= 32'b10010111010110010110100111110101;
12'b000010110011: dataA <= 32'b00000101101011001100110011110011;
12'b000010110100: dataA <= 32'b01000010111010100010100111101011;
12'b000010110101: dataA <= 32'b00000110011000001011101010110001;
12'b000010110110: dataA <= 32'b01100001001011110011001100010000;
12'b000010110111: dataA <= 32'b00001010101010000011001110101100;
12'b000010111000: dataA <= 32'b00011000111001101010000100000101;
12'b000010111001: dataA <= 32'b00000011010000101010011010001011;
12'b000010111010: dataA <= 32'b00110101010101010001100010000111;
12'b000010111011: dataA <= 32'b00001100100100010100110010111111;
12'b000010111100: dataA <= 32'b00110001000111010100101010010001;
12'b000010111101: dataA <= 32'b00000001110111101010101101110111;
12'b000010111110: dataA <= 32'b10011000001110100000010001100111;
12'b000010111111: dataA <= 32'b00001010001001110000001110001000;
12'b000011000000: dataA <= 32'b00010001011110001001110110100001;
12'b000011000001: dataA <= 32'b00001001001010001100110101000111;
12'b000011000010: dataA <= 32'b11011111010101111100001010001100;
12'b000011000011: dataA <= 32'b00001101000101000101001010100100;
12'b000011000100: dataA <= 32'b00000010111111110101001111001111;
12'b000011000101: dataA <= 32'b00001001001011101100100010001010;
12'b000011000110: dataA <= 32'b10011001100101001100011010001010;
12'b000011000111: dataA <= 32'b00000000101101000110011110000111;
12'b000011001000: dataA <= 32'b01101001010111000011000010010101;
12'b000011001001: dataA <= 32'b00001111001011011111000101110110;
12'b000011001010: dataA <= 32'b11100101111011110100011100110010;
12'b000011001011: dataA <= 32'b00001110110000101011001111100101;
12'b000011001100: dataA <= 32'b11010001110001100111101011001110;
12'b000011001101: dataA <= 32'b00001010000101011110011110111101;
12'b000011001110: dataA <= 32'b01101011001101111100111001110000;
12'b000011001111: dataA <= 32'b00000110011010011101010010101110;
12'b000011010000: dataA <= 32'b00011110010011011001100011001111;
12'b000011010001: dataA <= 32'b00001000111110100101011101011010;
12'b000011010010: dataA <= 32'b10001100111111100001110111101110;
12'b000011010011: dataA <= 32'b00001111010001011101100101111010;
12'b000011010100: dataA <= 32'b01010011010001011010000001001101;
12'b000011010101: dataA <= 32'b00001010110111011111100001110100;
12'b000011010110: dataA <= 32'b01101101001011110011111011101111;
12'b000011010111: dataA <= 32'b00001011101101011001000111011101;
12'b000011011000: dataA <= 32'b01101011000001011110101110001111;
12'b000011011001: dataA <= 32'b00001010000100001100011001011110;
12'b000011011010: dataA <= 32'b00011110000111001001001000100110;
12'b000011011011: dataA <= 32'b00001101001101001111010101011011;
12'b000011011100: dataA <= 32'b10100101001101010100100001110100;
12'b000011011101: dataA <= 32'b00000101001111001000111110110101;
12'b000011011110: dataA <= 32'b00101001010100111010101000100001;
12'b000011011111: dataA <= 32'b00001100010011011001100111001101;
12'b000011100000: dataA <= 32'b11100001101111001011101010001111;
12'b000011100001: dataA <= 32'b00001001100111010000110111001110;
12'b000011100010: dataA <= 32'b01010100011000100011100000101010;
12'b000011100011: dataA <= 32'b00001110010101011111010100110010;
12'b000011100100: dataA <= 32'b00101100100110100000010100101000;
12'b000011100101: dataA <= 32'b00001001110001011101001100011101;
12'b000011100110: dataA <= 32'b00100001011010110010000001101111;
12'b000011100111: dataA <= 32'b00001001001001100110000111100100;
12'b000011101000: dataA <= 32'b11011010100101100011100011110000;
12'b000011101001: dataA <= 32'b00000000101111000010110010011001;
12'b000011101010: dataA <= 32'b10101000111010101001001000000001;
12'b000011101011: dataA <= 32'b00000100111101100001000000110110;
12'b000011101100: dataA <= 32'b01001101001101110010010100101001;
12'b000011101101: dataA <= 32'b00000001101101010100010011101010;
12'b000011101110: dataA <= 32'b11001000101000111011100001001011;
12'b000011101111: dataA <= 32'b00001100010100011001011000001011;
12'b000011110000: dataA <= 32'b11100110001110001101000011011001;
12'b000011110001: dataA <= 32'b00000100110110100100111010000010;
12'b000011110010: dataA <= 32'b01000011000011110101000100011100;
12'b000011110011: dataA <= 32'b00001011101111100101000001000011;
12'b000011110100: dataA <= 32'b00001001010110110010010011010001;
12'b000011110101: dataA <= 32'b00001001001011010001000010011011;
12'b000011110110: dataA <= 32'b11100001001101010111010101011001;
12'b000011110111: dataA <= 32'b00001101011010101001101011110011;
12'b000011111000: dataA <= 32'b01100000000101101010000010101010;
12'b000011111001: dataA <= 32'b00000000101100101010000101011001;
12'b000011111010: dataA <= 32'b01001000011101010011001001000100;
12'b000011111011: dataA <= 32'b00001110010010010101100001010010;
12'b000011111100: dataA <= 32'b00100011001010000111101001011011;
12'b000011111101: dataA <= 32'b00001100001011100110110110101100;
12'b000011111110: dataA <= 32'b00011111100001110110101101110010;
12'b000011111111: dataA <= 32'b00001001100010011100010100111111;
12'b000100000000: dataA <= 32'b00000000000000110101010101010001;
12'b000100000001: dataA <= 32'b00000000000000000000000000000000;
12'b000100000010: dataA <= 32'b00001111100101111111100100111101;
12'b000100000011: dataA <= 32'b00001010101100010111010111100010;
12'b000100000100: dataA <= 32'b11000010101111101100101100110101;
12'b000100000101: dataA <= 32'b00001010100001011100001100011011;
12'b000100000110: dataA <= 32'b00101001111001111001110101001001;
12'b000100000111: dataA <= 32'b00001101000101100100100111000111;
12'b000100001000: dataA <= 32'b11011001011010100110011000010101;
12'b000100001001: dataA <= 32'b00000101001100001010111011110010;
12'b000100001010: dataA <= 32'b00000011000110011010010111101011;
12'b000100001011: dataA <= 32'b00000111011001010001110010100001;
12'b000100001100: dataA <= 32'b00100001001011101010011011101110;
12'b000100001101: dataA <= 32'b00001010001010000101011010101100;
12'b000100001110: dataA <= 32'b00011000111001100010000011000111;
12'b000100001111: dataA <= 32'b00000011010010100110010110001011;
12'b000100010000: dataA <= 32'b10110111001101001001110001101001;
12'b000100010001: dataA <= 32'b00001011100010010010110111010110;
12'b000100010010: dataA <= 32'b00110000111111010100001010010000;
12'b000100010011: dataA <= 32'b00000010111010101000101010000111;
12'b000100010100: dataA <= 32'b10010100010010001000010001001010;
12'b000100010101: dataA <= 32'b00001001001000101100001001111000;
12'b000100010110: dataA <= 32'b10010101100001111001110101000001;
12'b000100010111: dataA <= 32'b00001000101001001100111101011111;
12'b000100011000: dataA <= 32'b10100001010101111100001010001011;
12'b000100011001: dataA <= 32'b00001100000011000111010110100100;
12'b000100011010: dataA <= 32'b00000011001011110100011111001100;
12'b000100011011: dataA <= 32'b00001000101011101000011110000010;
12'b000100011100: dataA <= 32'b10011101101001010100101001101001;
12'b000100011101: dataA <= 32'b00000000110000000100101010011111;
12'b000100011110: dataA <= 32'b01101011010010111010110010110111;
12'b000100011111: dataA <= 32'b00001110101000011111000110000110;
12'b000100100000: dataA <= 32'b01101011111011110011101100110000;
12'b000100100001: dataA <= 32'b00001110001110101101001011110101;
12'b000100100010: dataA <= 32'b01010101111001111111101010101101;
12'b000100100011: dataA <= 32'b00001001000100011100011111000101;
12'b000100100100: dataA <= 32'b00101101001010000100111001101111;
12'b000100100101: dataA <= 32'b00000111011011011111010010110110;
12'b000100100110: dataA <= 32'b01011010010111001001000011010001;
12'b000100100111: dataA <= 32'b00001010011110101001011001010010;
12'b000100101000: dataA <= 32'b10001101000111010001010111001110;
12'b000100101001: dataA <= 32'b00001111001110011111100101110010;
12'b000100101010: dataA <= 32'b10010101010101010010010000110000;
12'b000100101011: dataA <= 32'b00001011010110100011011101111100;
12'b000100101100: dataA <= 32'b10101111000011110011001011101101;
12'b000100101101: dataA <= 32'b00001011101100011001001011100100;
12'b000100101110: dataA <= 32'b01101010111101101110111101101100;
12'b000100101111: dataA <= 32'b00001000100100001000100001101110;
12'b000100110000: dataA <= 32'b01011000001010111000101000000110;
12'b000100110001: dataA <= 32'b00001100101011010001011101011011;
12'b000100110010: dataA <= 32'b01100111001001011100110010010110;
12'b000100110011: dataA <= 32'b00000101010000001001000111000101;
12'b000100110100: dataA <= 32'b10101011010000110011000111000001;
12'b000100110101: dataA <= 32'b00001100110001011101101011001100;
12'b000100110110: dataA <= 32'b01100101101011000011001010001111;
12'b000100110111: dataA <= 32'b00001000100110010000111011011110;
12'b000100111000: dataA <= 32'b11010010011100100100000000101101;
12'b000100111001: dataA <= 32'b00001110110011100001010100101010;
12'b000100111010: dataA <= 32'b10101010011110010000010100001001;
12'b000100111011: dataA <= 32'b00001001110001011101001100100101;
12'b000100111100: dataA <= 32'b01100011011010100001110001110010;
12'b000100111101: dataA <= 32'b00001000001000100000000111100011;
12'b000100111110: dataA <= 32'b10011000100101100011100011110001;
12'b000100111111: dataA <= 32'b00000000110010000010111110001001;
12'b000101000000: dataA <= 32'b00101000110110010000110110100001;
12'b000101000001: dataA <= 32'b00000110011110100001000001001111;
12'b000101000010: dataA <= 32'b11001111010101101010100011101010;
12'b000101000011: dataA <= 32'b00000001110000010000010111100001;
12'b000101000100: dataA <= 32'b10000110110100111100000000101110;
12'b000101000101: dataA <= 32'b00001100010011011011011000001100;
12'b000101000110: dataA <= 32'b11100010001110010101000100011011;
12'b000101000111: dataA <= 32'b00000101011000100100111001111010;
12'b000101001000: dataA <= 32'b10000011001011110100010101111110;
12'b000101001001: dataA <= 32'b00001011101101100101000001000011;
12'b000101001010: dataA <= 32'b00001011011110101001110011110011;
12'b000101001011: dataA <= 32'b00001000101011010001001010011011;
12'b000101001100: dataA <= 32'b00100011001001101111100110011010;
12'b000101001101: dataA <= 32'b00001110011000101101100111110011;
12'b000101001110: dataA <= 32'b10011010000101011010010010101100;
12'b000101001111: dataA <= 32'b00000000101111100100000101001001;
12'b000101010000: dataA <= 32'b11000110100101001011011000000011;
12'b000101010001: dataA <= 32'b00001110001111011001100101001010;
12'b000101010010: dataA <= 32'b11100011001010010111101010011010;
12'b000101010011: dataA <= 32'b00001011101001100100110010101011;
12'b000101010100: dataA <= 32'b01100011011110001110101110010000;
12'b000101010101: dataA <= 32'b00001000000010011000010101010111;
12'b000101010110: dataA <= 32'b00000000000000111101100101010011;
12'b000101010111: dataA <= 32'b00000000000000000000000000000000;
12'b000101011000: dataA <= 32'b01010011101110010111100110011110;
12'b000101011001: dataA <= 32'b00001010001011011001011011010001;
12'b000101011010: dataA <= 32'b01000010110111110100001101010011;
12'b000101011011: dataA <= 32'b00001001000001010110001100100100;
12'b000101011100: dataA <= 32'b10101111110101101001110100101010;
12'b000101011101: dataA <= 32'b00001011100011100010100111010110;
12'b000101011110: dataA <= 32'b00011011011110101110001000110101;
12'b000101011111: dataA <= 32'b00000101001101001011000011101010;
12'b000101100000: dataA <= 32'b11000011010010010010000111001011;
12'b000101100001: dataA <= 32'b00001000011001010101111010010000;
12'b000101100010: dataA <= 32'b11100001001011100001111011101101;
12'b000101100011: dataA <= 32'b00001001001001000111100010101011;
12'b000101100100: dataA <= 32'b00011000111101011010010010001001;
12'b000101100101: dataA <= 32'b00000011110100100010010110000011;
12'b000101100110: dataA <= 32'b00111001000000111010010001001100;
12'b000101100111: dataA <= 32'b00001010000001010010111011100110;
12'b000101101000: dataA <= 32'b11110000110111010011101010001111;
12'b000101101001: dataA <= 32'b00000011111100100110100110011110;
12'b000101101010: dataA <= 32'b10001110010101110000010000101101;
12'b000101101011: dataA <= 32'b00001000101000100110000101100000;
12'b000101101100: dataA <= 32'b10010111100101101001110100000011;
12'b000101101101: dataA <= 32'b00001000001001001101000001101111;
12'b000101101110: dataA <= 32'b01100011010101111100001001101010;
12'b000101101111: dataA <= 32'b00001011000010001001011110101100;
12'b000101110000: dataA <= 32'b00000101010111110011101110101001;
12'b000101110001: dataA <= 32'b00001000001011100100011001110010;
12'b000101110010: dataA <= 32'b01100001101001010100111001001000;
12'b000101110011: dataA <= 32'b00000000110011000010110110110111;
12'b000101110100: dataA <= 32'b01101101001110110010010011011001;
12'b000101110101: dataA <= 32'b00001101100110100001000110010110;
12'b000101110110: dataA <= 32'b10101111110011110010111100101111;
12'b000101110111: dataA <= 32'b00001110001011101101000111110100;
12'b000101111000: dataA <= 32'b00011011111010010111101010101100;
12'b000101111001: dataA <= 32'b00001000000100011000011111001101;
12'b000101111010: dataA <= 32'b10101101000110001100111001101110;
12'b000101111011: dataA <= 32'b00001000111011100001010011000101;
12'b000101111100: dataA <= 32'b10010110010110111000100011110011;
12'b000101111101: dataA <= 32'b00001011111101101011010101001010;
12'b000101111110: dataA <= 32'b11001111001110111000110111001110;
12'b000101111111: dataA <= 32'b00001111001011100011100101101010;
12'b000110000000: dataA <= 32'b10010111011001001010100001010010;
12'b000110000001: dataA <= 32'b00001011110100100101011101111100;
12'b000110000010: dataA <= 32'b00101110111111101010011011001100;
12'b000110000011: dataA <= 32'b00001011001011011011001111100100;
12'b000110000100: dataA <= 32'b01101010111001111110111101001010;
12'b000110000101: dataA <= 32'b00000111100011000110101001111110;
12'b000110000110: dataA <= 32'b10010010001110100000010111000110;
12'b000110000111: dataA <= 32'b00001100001010010101100001010011;
12'b000110001000: dataA <= 32'b11100111000101100101000011011000;
12'b000110001001: dataA <= 32'b00000101010001001011001111000100;
12'b000110001010: dataA <= 32'b00101101001100101011100101100001;
12'b000110001011: dataA <= 32'b00001100101111100001101011001100;
12'b000110001100: dataA <= 32'b11101001101011000010101010001110;
12'b000110001101: dataA <= 32'b00000111100110010001000011101101;
12'b000110001110: dataA <= 32'b01001110100100100100100000110000;
12'b000110001111: dataA <= 32'b00001110110000100011010100101011;
12'b000110010000: dataA <= 32'b00100110011101111000010011101011;
12'b000110010001: dataA <= 32'b00001001110000011111001100110110;
12'b000110010010: dataA <= 32'b11100101011010010001100010010100;
12'b000110010011: dataA <= 32'b00000111101000011010000111011010;
12'b000110010100: dataA <= 32'b10010110101001100011110011110011;
12'b000110010101: dataA <= 32'b00000000110100000011001001111001;
12'b000110010110: dataA <= 32'b01100110110010000000110101000010;
12'b000110010111: dataA <= 32'b00000111111110100001000001011111;
12'b000110011000: dataA <= 32'b01010001011101100010100011101100;
12'b000110011001: dataA <= 32'b00000001110010001100011011010001;
12'b000110011010: dataA <= 32'b00000110111100111100100000110001;
12'b000110011011: dataA <= 32'b00001100110001011111011100001101;
12'b000110011100: dataA <= 32'b11011100001110011100110101011100;
12'b000110011101: dataA <= 32'b00000110011000100010110101110010;
12'b000110011110: dataA <= 32'b00000101010111110011100110111110;
12'b000110011111: dataA <= 32'b00001011001100100100111101000100;
12'b000110100000: dataA <= 32'b11001101100110011001110011110101;
12'b000110100001: dataA <= 32'b00001000001011010011001110010010;
12'b000110100010: dataA <= 32'b01100011001010000111100111011010;
12'b000110100011: dataA <= 32'b00001110110110101111011111101010;
12'b000110100100: dataA <= 32'b00010100001001010010100010001110;
12'b000110100101: dataA <= 32'b00000000110010011110000101000010;
12'b000110100110: dataA <= 32'b00000100110001001011100111000100;
12'b000110100111: dataA <= 32'b00001110001101011101101001000011;
12'b000110101000: dataA <= 32'b10100101000110101111011011011001;
12'b000110101001: dataA <= 32'b00001011001000100010110010101011;
12'b000110101010: dataA <= 32'b10100101011110011110101101101110;
12'b000110101011: dataA <= 32'b00000110100010010100011001101111;
12'b000110101100: dataA <= 32'b00000000000001001110000101110100;
12'b000110101101: dataA <= 32'b00000000000000000000000000000000;
12'b000110101110: dataA <= 32'b11010111110010101111100111111110;
12'b000110101111: dataA <= 32'b00001001101011011011011011000000;
12'b000110110000: dataA <= 32'b00000011000011101011011101010001;
12'b000110110001: dataA <= 32'b00000111100001010010010000100101;
12'b000110110010: dataA <= 32'b11110011101101100010000100001011;
12'b000110110011: dataA <= 32'b00001010100001100000100111100101;
12'b000110110100: dataA <= 32'b10011111011110111101111001010101;
12'b000110110101: dataA <= 32'b00000100101110001011001011011001;
12'b000110110110: dataA <= 32'b11000101011110000010000110101100;
12'b000110110111: dataA <= 32'b00001000111001011011111001111000;
12'b000110111000: dataA <= 32'b10100011000111010001011011001011;
12'b000110111001: dataA <= 32'b00001000101000001011101010101011;
12'b000110111010: dataA <= 32'b00011001000001001010100001101011;
12'b000110111011: dataA <= 32'b00000100010110011100010101111011;
12'b000110111100: dataA <= 32'b10111000111000110010100000101111;
12'b000110111101: dataA <= 32'b00001000100001010010111111101101;
12'b000110111110: dataA <= 32'b10101110110011001011001010001110;
12'b000110111111: dataA <= 32'b00000100111101100100100110101110;
12'b000111000000: dataA <= 32'b11001010011101011000010000110000;
12'b000111000001: dataA <= 32'b00000111100111100000000101010000;
12'b000111000010: dataA <= 32'b10011011101001100010000010100101;
12'b000111000011: dataA <= 32'b00000111001001001101001010000111;
12'b000111000100: dataA <= 32'b00100101010101111100001000101010;
12'b000111000101: dataA <= 32'b00001001100001001101100110101100;
12'b000111000110: dataA <= 32'b00000111100011110010111110000111;
12'b000111000111: dataA <= 32'b00000111101011100000011001101010;
12'b000111001000: dataA <= 32'b00100101101001011101001000001000;
12'b000111001001: dataA <= 32'b00000001010110000011000011000111;
12'b000111001010: dataA <= 32'b01101101001010101010000100011010;
12'b000111001011: dataA <= 32'b00001100100100100001000110100110;
12'b000111001100: dataA <= 32'b11110101101011101010001100101101;
12'b000111001101: dataA <= 32'b00001101101001101101000011110011;
12'b000111001110: dataA <= 32'b10100001111010101111101010001011;
12'b000111001111: dataA <= 32'b00000111000100010100100011010100;
12'b000111010000: dataA <= 32'b01101101000010001100111001101110;
12'b000111010001: dataA <= 32'b00001001111010100011010011001101;
12'b000111010010: dataA <= 32'b11010010011010100000010011110100;
12'b000111010011: dataA <= 32'b00001100111011101101010001000010;
12'b000111010100: dataA <= 32'b11001111010010101000010111001111;
12'b000111010101: dataA <= 32'b00001110101000100111100001100010;
12'b000111010110: dataA <= 32'b10011011011101000010110001010101;
12'b000111010111: dataA <= 32'b00001100010011101001011001111100;
12'b000111011000: dataA <= 32'b01101100110111100001111010101011;
12'b000111011001: dataA <= 32'b00001010101001011101001111100011;
12'b000111011010: dataA <= 32'b01101010110110001110111100101000;
12'b000111011011: dataA <= 32'b00000110100100000100110110001110;
12'b000111011100: dataA <= 32'b11001110010010001000010110000111;
12'b000111011101: dataA <= 32'b00001011101000011001100101010011;
12'b000111011110: dataA <= 32'b01100111000101101101010100011010;
12'b000111011111: dataA <= 32'b00000101010010001011010111001100;
12'b000111100000: dataA <= 32'b10101101001000101100000100100010;
12'b000111100001: dataA <= 32'b00001100101110100101101011001011;
12'b000111100010: dataA <= 32'b00101101100110110010011001101101;
12'b000111100011: dataA <= 32'b00000111000110010001000111110101;
12'b000111100100: dataA <= 32'b11001100101000101101000000110011;
12'b000111100101: dataA <= 32'b00001110101110100101010100100011;
12'b000111100110: dataA <= 32'b10100010011001100000010011001101;
12'b000111100111: dataA <= 32'b00001001101111100001001101000110;
12'b000111101000: dataA <= 32'b01100111010110000001100010110110;
12'b000111101001: dataA <= 32'b00000110101001010100001011010010;
12'b000111101010: dataA <= 32'b10010100101101100100000100010101;
12'b000111101011: dataA <= 32'b00000001110111000011010101110001;
12'b000111101100: dataA <= 32'b01100110110001101000110011100011;
12'b000111101101: dataA <= 32'b00001001011110100001000001110111;
12'b000111101110: dataA <= 32'b11010101100001011010110011001110;
12'b000111101111: dataA <= 32'b00000010010101001010100010111000;
12'b000111110000: dataA <= 32'b11000111001001000100110001010100;
12'b000111110001: dataA <= 32'b00001100101111100001011100011101;
12'b000111110010: dataA <= 32'b11011000001110011100110110111101;
12'b000111110011: dataA <= 32'b00000111011001100010110101101010;
12'b000111110100: dataA <= 32'b01000111100011110010111000011110;
12'b000111110101: dataA <= 32'b00001010101011100100111101000100;
12'b000111110110: dataA <= 32'b11010001101010001001100100110110;
12'b000111110111: dataA <= 32'b00000111101011010101010010001010;
12'b000111111000: dataA <= 32'b11100101001010011111101000111010;
12'b000111111001: dataA <= 32'b00001111010011110011011011100001;
12'b000111111010: dataA <= 32'b01001110001101001010110010010000;
12'b000111111011: dataA <= 32'b00000001010101011000000100110010;
12'b000111111100: dataA <= 32'b01000010111101001011110101100100;
12'b000111111101: dataA <= 32'b00001101101010100001101001000011;
12'b000111111110: dataA <= 32'b01100101000111000111001100010111;
12'b000111111111: dataA <= 32'b00001010000111100010110010101011;
12'b001000000000: dataA <= 32'b10101001011010101110011101101011;
12'b001000000001: dataA <= 32'b00000101100011010010011101111111;
12'b001000000010: dataA <= 32'b00000000000001010110010110010100;
12'b001000000011: dataA <= 32'b00000000000000000000000000000000;
12'b001000000100: dataA <= 32'b10011101110110111111001001011110;
12'b001000000101: dataA <= 32'b00001001001010011101011010110000;
12'b001000000110: dataA <= 32'b10000011001111101010101101001111;
12'b001000000111: dataA <= 32'b00000110000001001110011000101101;
12'b001000001000: dataA <= 32'b01110111100101010010010011101101;
12'b001000001001: dataA <= 32'b00001001000001011100100111110101;
12'b001000001010: dataA <= 32'b00100001011111000101011001110100;
12'b001000001011: dataA <= 32'b00000100110000001101010011001001;
12'b001000001100: dataA <= 32'b11001001100101111010000110001100;
12'b001000001101: dataA <= 32'b00001001111000100001111001101000;
12'b001000001110: dataA <= 32'b01100011000110111000111010101010;
12'b001000001111: dataA <= 32'b00001000001000010001110010100011;
12'b001000010000: dataA <= 32'b00011001000101000010110001001110;
12'b001000010001: dataA <= 32'b00000100110111011000010101110011;
12'b001000010010: dataA <= 32'b11110110110000101011000000110001;
12'b001000010011: dataA <= 32'b00000111000001010011000111110100;
12'b001000010100: dataA <= 32'b01101100101011001010101001101110;
12'b001000010101: dataA <= 32'b00000110011110100010100110111110;
12'b001000010110: dataA <= 32'b01001000100101000000100000110010;
12'b001000010111: dataA <= 32'b00000111001000011010000100111001;
12'b001000011000: dataA <= 32'b10011111101001010010010001100111;
12'b001000011001: dataA <= 32'b00000110101010001111010010011111;
12'b001000011010: dataA <= 32'b11100111010001111100001000001001;
12'b001000011011: dataA <= 32'b00001000000001010001101110101011;
12'b001000011100: dataA <= 32'b01001011101011101010001101000100;
12'b001000011101: dataA <= 32'b00000111001011011100011001011010;
12'b001000011110: dataA <= 32'b10101001100101100101010111101000;
12'b001000011111: dataA <= 32'b00000010011001000011001011011110;
12'b001000100000: dataA <= 32'b00101101000110011001110101111100;
12'b001000100001: dataA <= 32'b00001011100010100001000110101110;
12'b001000100010: dataA <= 32'b00111001100011011001101100001011;
12'b001000100011: dataA <= 32'b00001100100111101100111011110011;
12'b001000100100: dataA <= 32'b00100111111010111111001001101010;
12'b001000100101: dataA <= 32'b00000101100101010010100111010100;
12'b001000100110: dataA <= 32'b11101100111010010100101001001101;
12'b001000100111: dataA <= 32'b00001010111001100011001111010100;
12'b001000101000: dataA <= 32'b01001110100010001000010100010110;
12'b001000101001: dataA <= 32'b00001101111001101111001100111011;
12'b001000101010: dataA <= 32'b00010001011010010000010111001111;
12'b001000101011: dataA <= 32'b00001101100110101001011101011011;
12'b001000101100: dataA <= 32'b10011101011100111011010010010111;
12'b001000101101: dataA <= 32'b00001100010001101011010110000100;
12'b001000101110: dataA <= 32'b11101100110011010001001010001010;
12'b001000101111: dataA <= 32'b00001010001000011101001111011010;
12'b001000110000: dataA <= 32'b01101000110010100110101011100110;
12'b001000110001: dataA <= 32'b00000101000101000101000010011110;
12'b001000110010: dataA <= 32'b00001010011001110000010101101000;
12'b001000110011: dataA <= 32'b00001010100111011101100101010100;
12'b001000110100: dataA <= 32'b11101001000001110101010101011011;
12'b001000110101: dataA <= 32'b00000101110011001111011111001011;
12'b001000110110: dataA <= 32'b00101101000100101100100011000100;
12'b001000110111: dataA <= 32'b00001100001100101001100111001011;
12'b001000111000: dataA <= 32'b01110001011110101010001001101100;
12'b001000111001: dataA <= 32'b00000110000111010001001111110100;
12'b001000111010: dataA <= 32'b01001010110000110101100001010110;
12'b001000111011: dataA <= 32'b00001110001011100111010000100100;
12'b001000111100: dataA <= 32'b11011110011001001000100010101111;
12'b001000111101: dataA <= 32'b00001001101110100011001101010110;
12'b001000111110: dataA <= 32'b11101001010001110001100011111000;
12'b001000111111: dataA <= 32'b00000110001001001110001111000001;
12'b001001000000: dataA <= 32'b11010010110101100100010100110110;
12'b001001000001: dataA <= 32'b00000010011001000111011101100001;
12'b001001000010: dataA <= 32'b01100100101101011001000010100101;
12'b001001000011: dataA <= 32'b00001010111110100001000010001111;
12'b001001000100: dataA <= 32'b01011001100101010011000011010000;
12'b001001000101: dataA <= 32'b00000010110111000110101110101000;
12'b001001000110: dataA <= 32'b01001001010001001101010001110110;
12'b001001000111: dataA <= 32'b00001100101101100101011000100110;
12'b001001001000: dataA <= 32'b11010100010010100100101000011101;
12'b001001001001: dataA <= 32'b00001000011001100000110101101010;
12'b001001001010: dataA <= 32'b11001011101011101010001001111110;
12'b001001001011: dataA <= 32'b00001010001010100100111001000100;
12'b001001001100: dataA <= 32'b10010111110001111001100101010111;
12'b001001001101: dataA <= 32'b00000111001011010111010110000010;
12'b001001001110: dataA <= 32'b00100101000110101111011001111010;
12'b001001001111: dataA <= 32'b00001111010000110101010011010001;
12'b001001010000: dataA <= 32'b11001010010101000011000010010010;
12'b001001010001: dataA <= 32'b00000001111000010010001000101010;
12'b001001010010: dataA <= 32'b11000011000101001100010100100101;
12'b001001010011: dataA <= 32'b00001101001000100101101000111011;
12'b001001010100: dataA <= 32'b00100101000011010110101100110110;
12'b001001010101: dataA <= 32'b00001001000110100000101110100011;
12'b001001010110: dataA <= 32'b10101011010110110110001101001001;
12'b001001010111: dataA <= 32'b00000100100100001110100110010111;
12'b001001011000: dataA <= 32'b00000000000001100110100110110101;
12'b001001011001: dataA <= 32'b00000000000000000000000000000000;
12'b001001011010: dataA <= 32'b01100001110111010110101010011110;
12'b001001011011: dataA <= 32'b00001000101010100001011110011000;
12'b001001011100: dataA <= 32'b00000101011011011010001101001100;
12'b001001011101: dataA <= 32'b00000100100010001010011100111110;
12'b001001011110: dataA <= 32'b10111011011001001010100011101111;
12'b001001011111: dataA <= 32'b00000111100001011010100111110100;
12'b001001100000: dataA <= 32'b10100101011111001100111010010011;
12'b001001100001: dataA <= 32'b00000100110001001111011010110000;
12'b001001100010: dataA <= 32'b00001101101101101010000110001101;
12'b001001100011: dataA <= 32'b00001010110111100111111001011001;
12'b001001100100: dataA <= 32'b00100011000110101000011010001001;
12'b001001100101: dataA <= 32'b00000111001000010101111010100011;
12'b001001100110: dataA <= 32'b00011001000101000011010001010000;
12'b001001100111: dataA <= 32'b00000101111000010100011001110011;
12'b001001101000: dataA <= 32'b00110100101000101011100001010100;
12'b001001101001: dataA <= 32'b00000101100001010011001011110100;
12'b001001101010: dataA <= 32'b11101010100110111010001001101101;
12'b001001101011: dataA <= 32'b00000111111110011110100011001101;
12'b001001101100: dataA <= 32'b10000110101100110001000001010101;
12'b001001101101: dataA <= 32'b00000110001000010110000100101001;
12'b001001101110: dataA <= 32'b01100101101001001010100001001001;
12'b001001101111: dataA <= 32'b00000110001010010001011010110111;
12'b001001110000: dataA <= 32'b10101001001101111100000111101001;
12'b001001110001: dataA <= 32'b00000110100001010101110010101011;
12'b001001110010: dataA <= 32'b10001111110011011001101011100011;
12'b001001110011: dataA <= 32'b00000110101011011000011001010010;
12'b001001110100: dataA <= 32'b11101101100001101101010110101000;
12'b001001110101: dataA <= 32'b00000010111011000101010111100101;
12'b001001110110: dataA <= 32'b10101110111110001001110110111100;
12'b001001110111: dataA <= 32'b00001010000001100001000110111101;
12'b001001111000: dataA <= 32'b01111011011011001001001011101001;
12'b001001111001: dataA <= 32'b00001100000101101100110111101010;
12'b001001111010: dataA <= 32'b01101101110111010110101001001010;
12'b001001111011: dataA <= 32'b00000100100110010000101111010011;
12'b001001111100: dataA <= 32'b01101100110110010100101001001101;
12'b001001111101: dataA <= 32'b00001011111000100101001111010100;
12'b001001111110: dataA <= 32'b11001100101001110000010101010111;
12'b001001111111: dataA <= 32'b00001110110110101111000100111011;
12'b001010000000: dataA <= 32'b01010101011101111000010111001111;
12'b001010000001: dataA <= 32'b00001100100100101101011001011011;
12'b001010000010: dataA <= 32'b10100001100000111011110010111010;
12'b001010000011: dataA <= 32'b00001100101111101101010010000100;
12'b001010000100: dataA <= 32'b01101010101110111000111001101001;
12'b001010000101: dataA <= 32'b00001001001000011111001111010010;
12'b001010000110: dataA <= 32'b00100110101110110110011011000101;
12'b001010000111: dataA <= 32'b00000100000110000101001010101110;
12'b001010001000: dataA <= 32'b01000110100001011000010100101001;
12'b001010001001: dataA <= 32'b00001001100110100001101001010100;
12'b001010001010: dataA <= 32'b01101000111101111101010110011100;
12'b001010001011: dataA <= 32'b00000110010100010011100111001011;
12'b001010001100: dataA <= 32'b10101110111100110101000010000110;
12'b001010001101: dataA <= 32'b00001011101010101101100011000010;
12'b001010001110: dataA <= 32'b10110011010110011001111001001100;
12'b001010001111: dataA <= 32'b00000101001000010011010011110011;
12'b001010010000: dataA <= 32'b11001010111001000110000001111000;
12'b001010010001: dataA <= 32'b00001101101001101001001100101100;
12'b001010010010: dataA <= 32'b00011010011000111001000010110001;
12'b001010010011: dataA <= 32'b00001001101110100011001101100111;
12'b001010010100: dataA <= 32'b01101011001101100001100100011010;
12'b001010010101: dataA <= 32'b00000101101010001010010110111001;
12'b001010010110: dataA <= 32'b00010010111001100100010101110111;
12'b001010010111: dataA <= 32'b00000011011011001011101001010010;
12'b001010011000: dataA <= 32'b01100010101101001001010001100111;
12'b001010011001: dataA <= 32'b00001011111100100001000010011111;
12'b001010011010: dataA <= 32'b01011101100101010011010011010010;
12'b001010011011: dataA <= 32'b00000011111001000110110110010000;
12'b001010011100: dataA <= 32'b11001011011001010101100010111000;
12'b001010011101: dataA <= 32'b00001100001011100111011000110110;
12'b001010011110: dataA <= 32'b00001110011010100100011001011101;
12'b001010011111: dataA <= 32'b00001001011001100000110101100011;
12'b001010100000: dataA <= 32'b00001111110011011001101011011101;
12'b001010100001: dataA <= 32'b00001001101001100100111001001101;
12'b001010100010: dataA <= 32'b10011011110001101001100110011000;
12'b001010100011: dataA <= 32'b00000110101011011001011001111010;
12'b001010100100: dataA <= 32'b11100101000111000111001010111001;
12'b001010100101: dataA <= 32'b00001111001101110101001010111000;
12'b001010100110: dataA <= 32'b01000110011101000011100010110100;
12'b001010100111: dataA <= 32'b00000010111010001110001100101011;
12'b001010101000: dataA <= 32'b01000101010001001100100011100111;
12'b001010101001: dataA <= 32'b00001100000110101001100100111100;
12'b001010101010: dataA <= 32'b11100101000011100110001101010100;
12'b001010101011: dataA <= 32'b00001000000110011110101110011010;
12'b001010101100: dataA <= 32'b01101101010011000101101100000111;
12'b001010101101: dataA <= 32'b00000011000110001100101110101111;
12'b001010101110: dataA <= 32'b00000000000001110110100111010101;
12'b001010101111: dataA <= 32'b00000000000000000000000000000000;
12'b001010110000: dataA <= 32'b00111010111111010001011111001011;
12'b001010110001: dataA <= 32'b00000101001110101110111100001011;
12'b001010110010: dataA <= 32'b00101101110101000001000110000101;
12'b001010110011: dataA <= 32'b00000001010110001111101011000110;
12'b001010110100: dataA <= 32'b01101100001001010101100111111000;
12'b001010110101: dataA <= 32'b00000000110000010011001010010000;
12'b001010110110: dataA <= 32'b01101110110110011001101001101011;
12'b001010110111: dataA <= 32'b00001000110110101101100000010010;
12'b001010111000: dataA <= 32'b00110111100101000100100110110011;
12'b001010111001: dataA <= 32'b00001011101010111100110000100101;
12'b001010111010: dataA <= 32'b11100010111000001010100100101011;
12'b001010111011: dataA <= 32'b00000100010001111101010101100010;
12'b001010111100: dataA <= 32'b01100011001101101101111000011101;
12'b001010111101: dataA <= 32'b00001100010100001101010101100100;
12'b001010111110: dataA <= 32'b01010100010101110110101010011101;
12'b001010111111: dataA <= 32'b00000000110100100101011010000000;
12'b001011000000: dataA <= 32'b10010010101001000010000110101100;
12'b001011000001: dataA <= 32'b00001111010000010001000010111001;
12'b001011000010: dataA <= 32'b10010111110000100110011010111101;
12'b001011000011: dataA <= 32'b00000100010011000011010000110110;
12'b001011000100: dataA <= 32'b01110100110101010101100100111101;
12'b001011000101: dataA <= 32'b00000101010011101101011111101010;
12'b001011000110: dataA <= 32'b10100110101110000100000100110000;
12'b001011000111: dataA <= 32'b00000000110010111001010101110010;
12'b001011001000: dataA <= 32'b01111001100000110001000001101000;
12'b001011001001: dataA <= 32'b00000101110010001101001101010101;
12'b001011001010: dataA <= 32'b11110000100110101100100100010010;
12'b001011001011: dataA <= 32'b00001101111010101011110110111000;
12'b001011001100: dataA <= 32'b00011110100000111011101110010010;
12'b001011001101: dataA <= 32'b00000000101011100010111110110010;
12'b001011001110: dataA <= 32'b10101100001000100001100100101000;
12'b001011001111: dataA <= 32'b00000010100111011010100101001000;
12'b001011010000: dataA <= 32'b01111010100111010001010101001101;
12'b001011010001: dataA <= 32'b00000011010110010111011101101001;
12'b001011010010: dataA <= 32'b01011010100110010011010110101101;
12'b001011010011: dataA <= 32'b00001100001000100110110110001001;
12'b001011010100: dataA <= 32'b00010101100100001100011011110101;
12'b001011010101: dataA <= 32'b00001011000010100010100001111110;
12'b001011010110: dataA <= 32'b00101111010100001100000111110001;
12'b001011010111: dataA <= 32'b00000010000110101100100101101101;
12'b001011011000: dataA <= 32'b11110000111101111110001101011010;
12'b001011011001: dataA <= 32'b00000111100110101000100110010011;
12'b001011011010: dataA <= 32'b01010110101000011010000100101100;
12'b001011011011: dataA <= 32'b00000100001101100111000001001001;
12'b001011011100: dataA <= 32'b10010110110011001010010010101001;
12'b001011011101: dataA <= 32'b00000011010111100101110111000010;
12'b001011011110: dataA <= 32'b01010001110000001101000100110110;
12'b001011011111: dataA <= 32'b00000011001100110100111110001101;
12'b001011100000: dataA <= 32'b10011110101110101100001110010011;
12'b001011100001: dataA <= 32'b00001010010011110011011001101001;
12'b001011100010: dataA <= 32'b11011110100010100110010011011011;
12'b001011100011: dataA <= 32'b00000101001000110000100101010001;
12'b001011100100: dataA <= 32'b01101010011000111011000110001101;
12'b001011100101: dataA <= 32'b00000100010101101001011001110000;
12'b001011100110: dataA <= 32'b10011101101011000101111100011100;
12'b001011100111: dataA <= 32'b00000100100100100110101110011110;
12'b001011101000: dataA <= 32'b11001101001000100110001000111010;
12'b001011101001: dataA <= 32'b00000111001100100110111011100100;
12'b001011101010: dataA <= 32'b00100110101000110100111101010111;
12'b001011101011: dataA <= 32'b00000101010100001011101000101010;
12'b001011101100: dataA <= 32'b01011101011010001100111011110100;
12'b001011101101: dataA <= 32'b00001101111001110101101001000101;
12'b001011101110: dataA <= 32'b00010110111000101101100011111100;
12'b001011101111: dataA <= 32'b00001110001000100000111111101011;
12'b001011110000: dataA <= 32'b01110011000101101101011001011001;
12'b001011110001: dataA <= 32'b00001100111000011011110000001011;
12'b001011110010: dataA <= 32'b01101101101010110101011100011010;
12'b001011110011: dataA <= 32'b00000101100111101100110011011110;
12'b001011110100: dataA <= 32'b11001101100010001010111110101101;
12'b001011110101: dataA <= 32'b00001100101101011010111101100100;
12'b001011110110: dataA <= 32'b10111001100000110001001110101001;
12'b001011110111: dataA <= 32'b00000100101100011100110110100101;
12'b001011111000: dataA <= 32'b00111001001000110100101100010011;
12'b001011111001: dataA <= 32'b00000101110010101101001101010100;
12'b001011111010: dataA <= 32'b00100010110111100001111100101010;
12'b001011111011: dataA <= 32'b00000110100001100100010100011010;
12'b001011111100: dataA <= 32'b10001111110001110101111010011010;
12'b001011111101: dataA <= 32'b00001101011010000111100001101110;
12'b001011111110: dataA <= 32'b00101001110110010101100011111000;
12'b001011111111: dataA <= 32'b00000011000111110010101110001110;
12'b001100000000: dataA <= 32'b00100000110111000000111010000101;
12'b001100000001: dataA <= 32'b00000011001111010111000001011011;
12'b001100000010: dataA <= 32'b10101000100110110001110011100111;
12'b001100000011: dataA <= 32'b00000011011001010111100111101010;
12'b001100000100: dataA <= 32'b00000000000011010100011010110001;
12'b001100000101: dataA <= 32'b00000000000000000000000000000000;
12'b001100000110: dataA <= 32'b01111011000111100010001111001101;
12'b001100000111: dataA <= 32'b00000101001101101101000100010010;
12'b001100001000: dataA <= 32'b10100111111001010000100111100101;
12'b001100001001: dataA <= 32'b00000000110011001101100010110110;
12'b001100001010: dataA <= 32'b01110010010001001101010110111000;
12'b001100001011: dataA <= 32'b00000000101101010011000110101000;
12'b001100001100: dataA <= 32'b10101110111110101001111010001100;
12'b001100001101: dataA <= 32'b00001000010110101001100100100001;
12'b001100001110: dataA <= 32'b10110011101101000100000110010011;
12'b001100001111: dataA <= 32'b00001100001100111100111100011100;
12'b001100010000: dataA <= 32'b11100010111000011010000101001010;
12'b001100010001: dataA <= 32'b00000100001111111001011101101010;
12'b001100010010: dataA <= 32'b01100011001101011101110111011101;
12'b001100010011: dataA <= 32'b00001011110110001011001101100100;
12'b001100010100: dataA <= 32'b01011000010001100110101000111110;
12'b001100010101: dataA <= 32'b00000000110001100011011010011000;
12'b001100010110: dataA <= 32'b00010100100101010001100111001100;
12'b001100010111: dataA <= 32'b00001111010011010010111011001010;
12'b001100011000: dataA <= 32'b00010011101100010101111001011110;
12'b001100011001: dataA <= 32'b00000100010001000011001000101110;
12'b001100011010: dataA <= 32'b00110101000001001101010011111100;
12'b001100011011: dataA <= 32'b00000101010010101001100011110011;
12'b001100011100: dataA <= 32'b10101000110010000100000100101111;
12'b001100011101: dataA <= 32'b00000000101111110111011101111010;
12'b001100011110: dataA <= 32'b00110101101001000000100010000101;
12'b001100011111: dataA <= 32'b00000101110001001101000101001101;
12'b001100100000: dataA <= 32'b00110010101110101100110100010000;
12'b001100100001: dataA <= 32'b00001100111011100101111011010001;
12'b001100100010: dataA <= 32'b10100010100100111011001110010100;
12'b001100100011: dataA <= 32'b00000001001000100010111111000010;
12'b001100100100: dataA <= 32'b01110000001100110001000101100111;
12'b001100100101: dataA <= 32'b00000011100110011100100101100000;
12'b001100100110: dataA <= 32'b01111100110011100010000101001100;
12'b001100100111: dataA <= 32'b00000010110100010011011010000001;
12'b001100101000: dataA <= 32'b01011100100110010011010110101101;
12'b001100101001: dataA <= 32'b00001100101010100110111010011001;
12'b001100101010: dataA <= 32'b00010001100000001011101011010111;
12'b001100101011: dataA <= 32'b00001100100100100110100001101110;
12'b001100101100: dataA <= 32'b00101101011100001011010111110001;
12'b001100101101: dataA <= 32'b00000011000100101110101101100101;
12'b001100101110: dataA <= 32'b11101111000101101110001011111011;
12'b001100101111: dataA <= 32'b00001000100111101010101010010011;
12'b001100110000: dataA <= 32'b00011000100100100001010101001011;
12'b001100110001: dataA <= 32'b00000100001011100111000101011001;
12'b001100110010: dataA <= 32'b00011000101111010010110011001000;
12'b001100110011: dataA <= 32'b00000010110101100001110111001011;
12'b001100110100: dataA <= 32'b01001101101000001100010100010100;
12'b001100110101: dataA <= 32'b00000011101010110011000110000101;
12'b001100110110: dataA <= 32'b10100000101110101100011101110101;
12'b001100110111: dataA <= 32'b00001001110100101111100001111001;
12'b001100111000: dataA <= 32'b10100010100110010110100010011001;
12'b001100111001: dataA <= 32'b00000110000111110010101101100001;
12'b001100111010: dataA <= 32'b01101110011101000010100110001100;
12'b001100111011: dataA <= 32'b00000011110011100111011110001000;
12'b001100111100: dataA <= 32'b11011001101010110110011011011101;
12'b001100111101: dataA <= 32'b00000101100011101000110010001110;
12'b001100111110: dataA <= 32'b01001101000000010101100111111010;
12'b001100111111: dataA <= 32'b00000111001100100110111011011101;
12'b001101000000: dataA <= 32'b11101000101100110100011100011000;
12'b001101000001: dataA <= 32'b00000100110011000111100000111001;
12'b001101000010: dataA <= 32'b11011011011010001100111011010110;
12'b001101000011: dataA <= 32'b00001100111011101111110000111100;
12'b001101000100: dataA <= 32'b10010110110100100101000010111010;
12'b001101000101: dataA <= 32'b00001111001010100000111111101011;
12'b001101000110: dataA <= 32'b10110011001101100101011000011001;
12'b001101000111: dataA <= 32'b00001011111010010111110000001010;
12'b001101001000: dataA <= 32'b11101001101110101101101011011100;
12'b001101001001: dataA <= 32'b00000110100110101100110111001110;
12'b001101001010: dataA <= 32'b10001001010110010010111110101111;
12'b001101001011: dataA <= 32'b00001100101111011010111101011100;
12'b001101001100: dataA <= 32'b11110101101001000000101111001100;
12'b001101001101: dataA <= 32'b00000101001011011100110110011101;
12'b001101001110: dataA <= 32'b11111001010000110100001011110101;
12'b001101001111: dataA <= 32'b00000101110001101011010001010011;
12'b001101010000: dataA <= 32'b01100010110111101010101101001100;
12'b001101010001: dataA <= 32'b00001000000001101000010100100001;
12'b001101010010: dataA <= 32'b10001011101001100101111001011011;
12'b001101010011: dataA <= 32'b00001100011100000101011001011110;
12'b001101010100: dataA <= 32'b00100011111010001101100010110110;
12'b001101010101: dataA <= 32'b00000100000101110100110101111110;
12'b001101010110: dataA <= 32'b11100000110111010001011011000110;
12'b001101010111: dataA <= 32'b00000011001101010110111101100010;
12'b001101011000: dataA <= 32'b01101010101011000010010100100101;
12'b001101011001: dataA <= 32'b00000010010110010011100011110011;
12'b001101011010: dataA <= 32'b00000000000011010100111010110010;
12'b001101011011: dataA <= 32'b00000000000000000000000000000000;
12'b001101011100: dataA <= 32'b11111001010011110010101111010000;
12'b001101011101: dataA <= 32'b00000101101100101101001000011001;
12'b001101011110: dataA <= 32'b11100001111001101000101000100101;
12'b001101011111: dataA <= 32'b00000000110000001001011010100110;
12'b001101100000: dataA <= 32'b11110110011001000100110101110111;
12'b001101100001: dataA <= 32'b00000000101010010010111110111000;
12'b001101100010: dataA <= 32'b00101111000010111010001010101101;
12'b001101100011: dataA <= 32'b00000111010110100101101000110001;
12'b001101100100: dataA <= 32'b00101111110101000011110110010010;
12'b001101100101: dataA <= 32'b00001100101110111101001000011100;
12'b001101100110: dataA <= 32'b10100010111000101001010101101001;
12'b001101100111: dataA <= 32'b00000100001110110101101001110010;
12'b001101101000: dataA <= 32'b00100001001101010101100101111100;
12'b001101101001: dataA <= 32'b00001011010111001011000101100100;
12'b001101101010: dataA <= 32'b10011100001101010110010111111110;
12'b001101101011: dataA <= 32'b00000000101110011111011010110000;
12'b001101101100: dataA <= 32'b10011000100001100001100111001011;
12'b001101101101: dataA <= 32'b00001110110110010010110111010010;
12'b001101101110: dataA <= 32'b01001111101000001101001000011110;
12'b001101101111: dataA <= 32'b00000011110000000010111100011101;
12'b001101110000: dataA <= 32'b11110101001001000100110010111010;
12'b001101110001: dataA <= 32'b00000100110001100101100111110011;
12'b001101110010: dataA <= 32'b10101010110110000100000101001110;
12'b001101110011: dataA <= 32'b00000000101100110011100110000010;
12'b001101110100: dataA <= 32'b10110001110001011000010011100011;
12'b001101110101: dataA <= 32'b00000101110000001100111101000100;
12'b001101110110: dataA <= 32'b11110100110110100101000100001111;
12'b001101110111: dataA <= 32'b00001011011101100001111011100001;
12'b001101111000: dataA <= 32'b11100100100101000010101101010111;
12'b001101111001: dataA <= 32'b00000010000110100010111111001010;
12'b001101111010: dataA <= 32'b01110100010101000000100110100110;
12'b001101111011: dataA <= 32'b00000100100100100000100101111000;
12'b001101111100: dataA <= 32'b01111100111111110010100101101011;
12'b001101111101: dataA <= 32'b00000010010001010001010110010001;
12'b001101111110: dataA <= 32'b10100000100110011011100111001100;
12'b001101111111: dataA <= 32'b00001101001100101000111010101001;
12'b001110000000: dataA <= 32'b11001101011000001010111010011000;
12'b001110000001: dataA <= 32'b00001101100110101000100101011101;
12'b001110000010: dataA <= 32'b11101001100000001010100111110001;
12'b001110000011: dataA <= 32'b00000100000010110000110001011100;
12'b001110000100: dataA <= 32'b00101111001001011101111010111101;
12'b001110000101: dataA <= 32'b00001001100111101100101110010100;
12'b001110000110: dataA <= 32'b11011010100100111000110101101010;
12'b001110000111: dataA <= 32'b00000100101010100111000101101000;
12'b001110001000: dataA <= 32'b10011010101011011011100100000110;
12'b001110001001: dataA <= 32'b00000010010010011011110111001011;
12'b001110001010: dataA <= 32'b01001001100000001011100011110011;
12'b001110001011: dataA <= 32'b00000100001000110011001101111101;
12'b001110001100: dataA <= 32'b10100010110010101100101101010111;
12'b001110001101: dataA <= 32'b00001001010101101011101010001001;
12'b001110001110: dataA <= 32'b10100100100110000110100001010110;
12'b001110001111: dataA <= 32'b00000111000110110100110101110001;
12'b001110010000: dataA <= 32'b01110010100101001010010110101100;
12'b001110010001: dataA <= 32'b00000011010001100011011110100000;
12'b001110010010: dataA <= 32'b11010101100110100110101001111110;
12'b001110010011: dataA <= 32'b00000111000010101010110101111110;
12'b001110010100: dataA <= 32'b11001100111000001100110110111001;
12'b001110010101: dataA <= 32'b00000111101100100110111111010101;
12'b001110010110: dataA <= 32'b01101010110000110011111011011010;
12'b001110010111: dataA <= 32'b00000100110010000101010101001001;
12'b001110011000: dataA <= 32'b01010111010110000100111010110111;
12'b001110011001: dataA <= 32'b00001011111100101011111000110100;
12'b001110011010: dataA <= 32'b01011000110000011100100001111000;
12'b001110011011: dataA <= 32'b00001111001101100000111111101100;
12'b001110011100: dataA <= 32'b00110001010101011101000111011001;
12'b001110011101: dataA <= 32'b00001010111011010001101000011010;
12'b001110011110: dataA <= 32'b00100101110010011101111010011101;
12'b001110011111: dataA <= 32'b00000111100110101110111110111111;
12'b001110100000: dataA <= 32'b10000111001110011011001110110010;
12'b001110100001: dataA <= 32'b00001100110001011010111001011100;
12'b001110100010: dataA <= 32'b11110001110001011000011111001111;
12'b001110100011: dataA <= 32'b00000101101010011110110110001101;
12'b001110100100: dataA <= 32'b10110101011100110011101011010110;
12'b001110100101: dataA <= 32'b00000101110000101001010101011011;
12'b001110100110: dataA <= 32'b11100100110111110011001101001110;
12'b001110100111: dataA <= 32'b00001001100001101100011000111000;
12'b001110101000: dataA <= 32'b01000111100001011101101000011011;
12'b001110101001: dataA <= 32'b00001010111101000011001101001110;
12'b001110101010: dataA <= 32'b11011111111001111101100010010100;
12'b001110101011: dataA <= 32'b00000101000100110100111101101101;
12'b001110101100: dataA <= 32'b10100010110111100001111011100111;
12'b001110101101: dataA <= 32'b00000011101011011000111001101010;
12'b001110101110: dataA <= 32'b00101100101111001010100101100100;
12'b001110101111: dataA <= 32'b00000001110100001111011011110100;
12'b001110110000: dataA <= 32'b00000000000011001101011010010011;
12'b001110110001: dataA <= 32'b00000000000000000000000000000000;
12'b001110110010: dataA <= 32'b01110111011011110011011111010011;
12'b001110110011: dataA <= 32'b00000101101011101101001100101001;
12'b001110110100: dataA <= 32'b11011011111010000000011001100101;
12'b001110110101: dataA <= 32'b00000000101101000111010010001110;
12'b001110110110: dataA <= 32'b01111010100000111100100101010110;
12'b001110110111: dataA <= 32'b00000001101000010010111011010001;
12'b001110111000: dataA <= 32'b10101111001011000010101010101110;
12'b001110111001: dataA <= 32'b00000110110101100001101001000000;
12'b001110111010: dataA <= 32'b01101001111001000011010101110001;
12'b001110111011: dataA <= 32'b00001100101111111101010100011011;
12'b001110111100: dataA <= 32'b10100100111100111000110110101000;
12'b001110111101: dataA <= 32'b00000100101101110001110001111010;
12'b001110111110: dataA <= 32'b11011111001101001101000100111011;
12'b001110111111: dataA <= 32'b00001010011000001010111001100011;
12'b001111000000: dataA <= 32'b11100000001101001110000110011101;
12'b001111000001: dataA <= 32'b00000000101011011101011011000000;
12'b001111000010: dataA <= 32'b00011010011101110001010111101011;
12'b001111000011: dataA <= 32'b00001110011000010010110011011011;
12'b001111000100: dataA <= 32'b11001011100000001100010110111110;
12'b001111000101: dataA <= 32'b00000100001110000010110000010100;
12'b001111000110: dataA <= 32'b10110011010000111100100001110111;
12'b001111000111: dataA <= 32'b00000100101111100001100111110100;
12'b001111001000: dataA <= 32'b10101010111010000100000101001100;
12'b001111001001: dataA <= 32'b00000001001001101111101110001010;
12'b001111001010: dataA <= 32'b01101011110101110000010100100010;
12'b001111001011: dataA <= 32'b00000101101111001100110101000100;
12'b001111001100: dataA <= 32'b01110100111110011101010100001101;
12'b001111001101: dataA <= 32'b00001001111110011011111011101010;
12'b001111001110: dataA <= 32'b01100110100101001010011100111001;
12'b001111001111: dataA <= 32'b00000011000100100010111111001011;
12'b001111010000: dataA <= 32'b01111000100001011000010111100110;
12'b001111010001: dataA <= 32'b00000101100011100010100110010000;
12'b001111010010: dataA <= 32'b10111101001011110011010110001010;
12'b001111010011: dataA <= 32'b00000010001111001111001110100001;
12'b001111010100: dataA <= 32'b11100010100110011011100111001100;
12'b001111010101: dataA <= 32'b00001101101110101000111110110001;
12'b001111010110: dataA <= 32'b10001011010000010010001001111000;
12'b001111010111: dataA <= 32'b00001110101000101010101001010101;
12'b001111011000: dataA <= 32'b10100111100000011010000111010001;
12'b001111011001: dataA <= 32'b00000101100001110010111001011100;
12'b001111011010: dataA <= 32'b00101101010001010101101001011101;
12'b001111011011: dataA <= 32'b00001010001000101110110110010100;
12'b001111011100: dataA <= 32'b11011110100001001000100110001001;
12'b001111011101: dataA <= 32'b00000101101001100111001010000000;
12'b001111011110: dataA <= 32'b00011100101011011100000101000101;
12'b001111011111: dataA <= 32'b00000001110000010101110011001100;
12'b001111100000: dataA <= 32'b01000111011000001010110011010001;
12'b001111100001: dataA <= 32'b00000101000111110001010101110101;
12'b001111100010: dataA <= 32'b11100010110010100100111100011001;
12'b001111100011: dataA <= 32'b00001000110101100111101010011001;
12'b001111100100: dataA <= 32'b10100110100101110110100000110100;
12'b001111100101: dataA <= 32'b00000111100110110100111110000001;
12'b001111100110: dataA <= 32'b10110100101101010001110111001011;
12'b001111100111: dataA <= 32'b00000011010000100001011110111000;
12'b001111101000: dataA <= 32'b10010011100010010110111000011110;
12'b001111101001: dataA <= 32'b00001000000010101010111001101110;
12'b001111101010: dataA <= 32'b01001110110000001100000101111000;
12'b001111101011: dataA <= 32'b00001000001100100111000011000110;
12'b001111101100: dataA <= 32'b00101100110100110011011010011011;
12'b001111101101: dataA <= 32'b00000100010000000011001001011001;
12'b001111101110: dataA <= 32'b00010101010001111100111001111000;
12'b001111101111: dataA <= 32'b00001010011110100101111000110100;
12'b001111110000: dataA <= 32'b00011000110000011011110001010101;
12'b001111110001: dataA <= 32'b00001111010000100000111111101101;
12'b001111110010: dataA <= 32'b01101111011101010100110110011000;
12'b001111110011: dataA <= 32'b00001001011100001101100100101001;
12'b001111110100: dataA <= 32'b10011111110010010110001000111110;
12'b001111110101: dataA <= 32'b00001000100110101111000010100111;
12'b001111110110: dataA <= 32'b01000111000110011011001110010101;
12'b001111110111: dataA <= 32'b00001100010011011010111001011100;
12'b001111111000: dataA <= 32'b11101011110101110000011111010010;
12'b001111111001: dataA <= 32'b00000110001001011110110110000101;
12'b001111111010: dataA <= 32'b01110011100100111011001010111000;
12'b001111111011: dataA <= 32'b00000101101111100111011001011011;
12'b001111111100: dataA <= 32'b10100100111011110011111101010001;
12'b001111111101: dataA <= 32'b00001011000010101110100001001000;
12'b001111111110: dataA <= 32'b11000101010101010101010111011011;
12'b001111111111: dataA <= 32'b00001001011110000011000001000101;
12'b010000000000: dataA <= 32'b11011001110101110101100010010001;
12'b010000000001: dataA <= 32'b00000110100011110101000101100101;
12'b010000000010: dataA <= 32'b10100010110111101010101100101001;
12'b010000000011: dataA <= 32'b00000100001001011000111001110010;
12'b010000000100: dataA <= 32'b10101110110111010011000111000100;
12'b010000000101: dataA <= 32'b00000001010010001101010111110100;
12'b010000000110: dataA <= 32'b00000000000011000101101010010100;
12'b010000000111: dataA <= 32'b00000000000000000000000000000000;
12'b010000001000: dataA <= 32'b11110011100011110100001110110110;
12'b010000001001: dataA <= 32'b00000110001010101011010001000000;
12'b010000001010: dataA <= 32'b00010111111010010000101010100110;
12'b010000001011: dataA <= 32'b00000000101010000111000101111111;
12'b010000001100: dataA <= 32'b11111100101100111100000100110101;
12'b010000001101: dataA <= 32'b00000010100101010010110111100001;
12'b010000001110: dataA <= 32'b01101101001111001010111010101111;
12'b010000001111: dataA <= 32'b00000110010101011101101001011000;
12'b010000010000: dataA <= 32'b11100011111001001011000101110000;
12'b010000010001: dataA <= 32'b00001100110001111001011100100010;
12'b010000010010: dataA <= 32'b10100100111101001000100111001000;
12'b010000010011: dataA <= 32'b00000101001011101101110110000010;
12'b010000010100: dataA <= 32'b10011101001101000100110011111001;
12'b010000010101: dataA <= 32'b00001001011001001010110001100011;
12'b010000010110: dataA <= 32'b01100110010000111101100100111100;
12'b010000010111: dataA <= 32'b00000001001000011011011011010001;
12'b010000011000: dataA <= 32'b11011110011110000001011000001011;
12'b010000011001: dataA <= 32'b00001101011010010100101111100011;
12'b010000011010: dataA <= 32'b00001001010100001011100101011101;
12'b010000011011: dataA <= 32'b00000100001101000100100100010100;
12'b010000011100: dataA <= 32'b00110001010100111100000000110101;
12'b010000011101: dataA <= 32'b00000100101110011111100111110101;
12'b010000011110: dataA <= 32'b11101010111110000100000101101011;
12'b010000011111: dataA <= 32'b00000001100111101011110010010010;
12'b010000100000: dataA <= 32'b11100101111010001000010110000001;
12'b010000100001: dataA <= 32'b00000101101110001110101101000011;
12'b010000100010: dataA <= 32'b00110101000110010101010100101100;
12'b010000100011: dataA <= 32'b00001000011110010101110111110011;
12'b010000100100: dataA <= 32'b11101000101001011010001011111010;
12'b010000100101: dataA <= 32'b00000100000010100011000011001011;
12'b010000100110: dataA <= 32'b01111100101001110000011000000110;
12'b010000100111: dataA <= 32'b00000111000011100100100110101000;
12'b010000101000: dataA <= 32'b11111101010111110100000110101010;
12'b010000101001: dataA <= 32'b00000010001101001111000110101001;
12'b010000101010: dataA <= 32'b01100100100110011011110111101100;
12'b010000101011: dataA <= 32'b00001101110001101001000011000010;
12'b010000101100: dataA <= 32'b01001011001000100001101000111001;
12'b010000101101: dataA <= 32'b00001111001011101100101101001101;
12'b010000101110: dataA <= 32'b01100011100100101001010111010001;
12'b010000101111: dataA <= 32'b00000111000001110011000001010100;
12'b010000110000: dataA <= 32'b00101011010101001101011000011110;
12'b010000110001: dataA <= 32'b00001011001001101110111010010100;
12'b010000110010: dataA <= 32'b11100000100001100000010110101000;
12'b010000110011: dataA <= 32'b00000110001000100101001110010000;
12'b010000110100: dataA <= 32'b10011110101011011100100110000100;
12'b010000110101: dataA <= 32'b00000010001110010001101111001100;
12'b010000110110: dataA <= 32'b00000101001100010010000011001111;
12'b010000110111: dataA <= 32'b00000101100110101111011101101101;
12'b010000111000: dataA <= 32'b11100100110010011101001011011011;
12'b010000111001: dataA <= 32'b00001000010101100011101110101001;
12'b010000111010: dataA <= 32'b10101000101001100110010000110001;
12'b010000111011: dataA <= 32'b00001000100110110101000110010001;
12'b010000111100: dataA <= 32'b00110100110101100001110111101011;
12'b010000111101: dataA <= 32'b00000011001110011101011111001001;
12'b010000111110: dataA <= 32'b10001111011010000110110110111110;
12'b010000111111: dataA <= 32'b00001001100010101010111101011110;
12'b010001000000: dataA <= 32'b11001110101000001011010100110111;
12'b010001000001: dataA <= 32'b00001000101100100111000110110110;
12'b010001000010: dataA <= 32'b11101100111000111010111001011100;
12'b010001000011: dataA <= 32'b00000100001111000010111101101000;
12'b010001000100: dataA <= 32'b10010011001101110100111000111000;
12'b010001000101: dataA <= 32'b00001001011110011111111000110011;
12'b010001000110: dataA <= 32'b10011010101100011011010000110010;
12'b010001000111: dataA <= 32'b00001111010011100000111111100101;
12'b010001001000: dataA <= 32'b11101011100001010100100101011000;
12'b010001001001: dataA <= 32'b00001000011100001011011100111000;
12'b010001001010: dataA <= 32'b10011011110010000110000111011110;
12'b010001001011: dataA <= 32'b00001001100111101101001010010111;
12'b010001001100: dataA <= 32'b00000110111010100011011101110111;
12'b010001001101: dataA <= 32'b00001100010101011100110101011100;
12'b010001001110: dataA <= 32'b11100101111010001000011111010100;
12'b010001001111: dataA <= 32'b00000110101000100000110101110101;
12'b010001010000: dataA <= 32'b00101111101000111010101001111000;
12'b010001010001: dataA <= 32'b00000101101110100101011101100011;
12'b010001010010: dataA <= 32'b01100100111011110100101101010011;
12'b010001010011: dataA <= 32'b00001100000011110010100101100000;
12'b010001010100: dataA <= 32'b10000011001001001101000110011010;
12'b010001010101: dataA <= 32'b00000111111110000010110100110101;
12'b010001010110: dataA <= 32'b10010011110001101101100001101111;
12'b010001010111: dataA <= 32'b00000111100011110011001101011101;
12'b010001011000: dataA <= 32'b10100100111011110011011101001011;
12'b010001011001: dataA <= 32'b00000100101000011000110101111010;
12'b010001011010: dataA <= 32'b01101110111011010011101000000011;
12'b010001011011: dataA <= 32'b00000001001111001011001111101101;
12'b010001011100: dataA <= 32'b00000000000010110110001001110101;
12'b010001011101: dataA <= 32'b00000000000000000000000000000000;
12'b010001011110: dataA <= 32'b01101111101011110100111110011000;
12'b010001011111: dataA <= 32'b00000111001010101001010101010000;
12'b010001100000: dataA <= 32'b11010001110010101000101011000111;
12'b010001100001: dataA <= 32'b00000001101000000100111101101110;
12'b010001100010: dataA <= 32'b01111100111000111011100100010100;
12'b010001100011: dataA <= 32'b00000011100011010100110011101010;
12'b010001100100: dataA <= 32'b01101011010011010011011010110000;
12'b010001100101: dataA <= 32'b00000101110100011001100101110000;
12'b010001100110: dataA <= 32'b01011101111001010010110101110000;
12'b010001100111: dataA <= 32'b00001100010011110101101000101010;
12'b010001101000: dataA <= 32'b10100100111101100000011000000111;
12'b010001101001: dataA <= 32'b00000101001010100111111010001010;
12'b010001101010: dataA <= 32'b10011101001101000100100010110111;
12'b010001101011: dataA <= 32'b00001000011001001100101001100011;
12'b010001101100: dataA <= 32'b00101010010100110101010011111011;
12'b010001101101: dataA <= 32'b00000010000110011001010111100010;
12'b010001101110: dataA <= 32'b01100010011110010001011000101011;
12'b010001101111: dataA <= 32'b00001011111100010110101011100100;
12'b010001110000: dataA <= 32'b10000111001100001010110011111100;
12'b010001110001: dataA <= 32'b00000100101011000110011100010011;
12'b010001110010: dataA <= 32'b11101111011100111011100000110010;
12'b010001110011: dataA <= 32'b00000101001101011011100111100101;
12'b010001110100: dataA <= 32'b11101011000010000100000110001011;
12'b010001110101: dataA <= 32'b00000010100101100101110110011010;
12'b010001110110: dataA <= 32'b10011111111010100000010111100001;
12'b010001110111: dataA <= 32'b00000101101101010000100101000011;
12'b010001111000: dataA <= 32'b11110011001110001101100101001011;
12'b010001111001: dataA <= 32'b00000110111110001111110011110011;
12'b010001111010: dataA <= 32'b01101010101101100001111010111011;
12'b010001111011: dataA <= 32'b00000101100001100011000011001100;
12'b010001111100: dataA <= 32'b11111100110110001000011001000110;
12'b010001111101: dataA <= 32'b00001000000010100110101010111000;
12'b010001111110: dataA <= 32'b00111001011111110100110111001001;
12'b010001111111: dataA <= 32'b00000010101011001111000010111010;
12'b010010000000: dataA <= 32'b10100110101010011100001000001100;
12'b010010000001: dataA <= 32'b00001101010011101001000111001010;
12'b010010000010: dataA <= 32'b00001001000000110001000111111001;
12'b010010000011: dataA <= 32'b00001111001110101110110101000101;
12'b010010000100: dataA <= 32'b00011111100100111000110111010000;
12'b010010000101: dataA <= 32'b00001000100001110011000101010100;
12'b010010000110: dataA <= 32'b01101001011001000101000110111101;
12'b010010000111: dataA <= 32'b00001011101010110001000010001100;
12'b010010001000: dataA <= 32'b00100100100101111000010111101000;
12'b010010001001: dataA <= 32'b00000110101000100011001110101001;
12'b010010001010: dataA <= 32'b00100000101011010101000111100011;
12'b010010001011: dataA <= 32'b00000010001011001101100111001101;
12'b010010001100: dataA <= 32'b00000011000000100001100011001110;
12'b010010001101: dataA <= 32'b00000110100101101011100001100101;
12'b010010001110: dataA <= 32'b01100110110110010101011010011100;
12'b010010001111: dataA <= 32'b00000111110101011111101110110010;
12'b010010010000: dataA <= 32'b10101010101101010110000000101110;
12'b010010010001: dataA <= 32'b00001001100111110011001110100001;
12'b010010010010: dataA <= 32'b10110110111101110001100111101011;
12'b010010010011: dataA <= 32'b00000011101100011011011111011001;
12'b010010010100: dataA <= 32'b01001101010101110110110101011110;
12'b010010010101: dataA <= 32'b00001010100011101011000001001110;
12'b010010010110: dataA <= 32'b00010010100100001010110100010110;
12'b010010010111: dataA <= 32'b00001000101100100111000110100111;
12'b010010011000: dataA <= 32'b11101100111101000010010111111100;
12'b010010011001: dataA <= 32'b00000100101101000010110010000000;
12'b010010011010: dataA <= 32'b00010011001001110100111000011000;
12'b010010011011: dataA <= 32'b00000111111110011001111000111011;
12'b010010011100: dataA <= 32'b01011100101100100010100000101111;
12'b010010011101: dataA <= 32'b00001110110110100000111111010110;
12'b010010011110: dataA <= 32'b10100111100101001100010100110110;
12'b010010011111: dataA <= 32'b00000110111100001001010101001000;
12'b010010100000: dataA <= 32'b10010101101101110110000101111101;
12'b010010100001: dataA <= 32'b00001010000111101101001101111111;
12'b010010100010: dataA <= 32'b11000110110010100011101100111001;
12'b010010100011: dataA <= 32'b00001011010110011100110101011011;
12'b010010100100: dataA <= 32'b11100001111010100000011110010111;
12'b010010100101: dataA <= 32'b00000111101000100000110101101101;
12'b010010100110: dataA <= 32'b00101011101101001010011000111001;
12'b010010100111: dataA <= 32'b00000101101101100001011101100011;
12'b010010101000: dataA <= 32'b01100110111111101101011100110101;
12'b010010101001: dataA <= 32'b00001101000101110100101101111000;
12'b010010101010: dataA <= 32'b00000010111101000100100101011010;
12'b010010101011: dataA <= 32'b00000110011110000010101000101101;
12'b010010101100: dataA <= 32'b01001111101101100101010010001101;
12'b010010101101: dataA <= 32'b00001001000011110001010101001101;
12'b010010101110: dataA <= 32'b10100100111011110011111101101101;
12'b010010101111: dataA <= 32'b00000101100111011010110010000010;
12'b010010110000: dataA <= 32'b00110001000011010100011001000100;
12'b010010110001: dataA <= 32'b00000001001100001011000111100110;
12'b010010110010: dataA <= 32'b00000000000010101110011000110101;
12'b010010110011: dataA <= 32'b00000000000000000000000000000000;
12'b010010110100: dataA <= 32'b01101011101111101101101101011011;
12'b010010110101: dataA <= 32'b00000111101001100101011001101000;
12'b010010110110: dataA <= 32'b10001101101110111001001100001001;
12'b010010110111: dataA <= 32'b00000010000101000110110001010110;
12'b010010111000: dataA <= 32'b00111101000100111011010011110010;
12'b010010111001: dataA <= 32'b00000100100010010110101111110011;
12'b010010111010: dataA <= 32'b01101001010111010011111010110001;
12'b010010111011: dataA <= 32'b00000101010011010101100110001000;
12'b010010111100: dataA <= 32'b11010111111001011010100101101111;
12'b010010111101: dataA <= 32'b00001011110100110001110000111001;
12'b010010111110: dataA <= 32'b11100101000001111000011000101000;
12'b010010111111: dataA <= 32'b00000110001001100001111010010010;
12'b010011000000: dataA <= 32'b01011011001000111100000010010101;
12'b010011000001: dataA <= 32'b00000111011001001110100101101011;
12'b010011000010: dataA <= 32'b10101110011000101100110010111001;
12'b010011000011: dataA <= 32'b00000011000100010111010011110010;
12'b010011000100: dataA <= 32'b11100100011110100001101000101100;
12'b010011000101: dataA <= 32'b00001010111110011010100111011100;
12'b010011000110: dataA <= 32'b11000101000000010010000010111010;
12'b010011000111: dataA <= 32'b00000101001010001010010000011010;
12'b010011001000: dataA <= 32'b01101011100000111011010000101111;
12'b010011001001: dataA <= 32'b00000101001100010111100011011110;
12'b010011001010: dataA <= 32'b00101011000110000100000110101010;
12'b010011001011: dataA <= 32'b00000100000011011111110110100011;
12'b010011001100: dataA <= 32'b00011011111010111000101001000001;
12'b010011001101: dataA <= 32'b00000101101101010010100001000011;
12'b010011001110: dataA <= 32'b10110011010101111101100101101010;
12'b010011001111: dataA <= 32'b00000101111110001011101011110100;
12'b010011010000: dataA <= 32'b11101100110101110001111001011100;
12'b010011010001: dataA <= 32'b00000111000001100011000011001100;
12'b010011010010: dataA <= 32'b00111101000010100000011010000111;
12'b010011010011: dataA <= 32'b00001001100011101000101111010001;
12'b010011010100: dataA <= 32'b10110111101011101101101000001001;
12'b010011010101: dataA <= 32'b00000011001001001110111011000010;
12'b010011010110: dataA <= 32'b00101000101110011100011000101100;
12'b010011010111: dataA <= 32'b00001100110101100111000111010011;
12'b010011011000: dataA <= 32'b10001000111001000000100110111001;
12'b010011011001: dataA <= 32'b00001111010001101110111000111100;
12'b010011011010: dataA <= 32'b11011011100101001000100111010000;
12'b010011011011: dataA <= 32'b00001010000001110001001101010011;
12'b010011011100: dataA <= 32'b01100111011100111100100101011101;
12'b010011011101: dataA <= 32'b00001100001100101111000110001100;
12'b010011011110: dataA <= 32'b01100110100110010000011000001000;
12'b010011011111: dataA <= 32'b00000111100111100011001110111001;
12'b010011100000: dataA <= 32'b01100010101011001101101000100100;
12'b010011100001: dataA <= 32'b00000010101001001001011111000101;
12'b010011100010: dataA <= 32'b11000010111000110001000011101100;
12'b010011100011: dataA <= 32'b00000111100101100111100101011100;
12'b010011100100: dataA <= 32'b10100110110110001101011000111101;
12'b010011100101: dataA <= 32'b00000111010101011011101110111010;
12'b010011100110: dataA <= 32'b11101100110101000101110000101011;
12'b010011100111: dataA <= 32'b00001010001000110011010110101001;
12'b010011101000: dataA <= 32'b00110111000110000001101000001011;
12'b010011101001: dataA <= 32'b00000100001011010111011011101010;
12'b010011101010: dataA <= 32'b11001011001101011110100100011100;
12'b010011101011: dataA <= 32'b00001100000101101011000100111101;
12'b010011101100: dataA <= 32'b01010100100000011010000011110100;
12'b010011101101: dataA <= 32'b00001001001101100101001010001111;
12'b010011101110: dataA <= 32'b11101101000101001010000110111100;
12'b010011101111: dataA <= 32'b00000100101100000100101010010000;
12'b010011110000: dataA <= 32'b11010011000101101100100111011000;
12'b010011110001: dataA <= 32'b00000110011110010011110101000010;
12'b010011110010: dataA <= 32'b10011110101000101010000000101101;
12'b010011110011: dataA <= 32'b00001110011000100000111111000110;
12'b010011110100: dataA <= 32'b01100011100101001011110100010101;
12'b010011110101: dataA <= 32'b00000101111011000111001001100000;
12'b010011110110: dataA <= 32'b10010001101001101110000100111100;
12'b010011110111: dataA <= 32'b00001011001000101011010001100111;
12'b010011111000: dataA <= 32'b10001000101010101011111011111011;
12'b010011111001: dataA <= 32'b00001010110111011110110101011011;
12'b010011111010: dataA <= 32'b10011011111010111000101101111001;
12'b010011111011: dataA <= 32'b00001000001000100010110101011101;
12'b010011111100: dataA <= 32'b11100101110001010010000111111001;
12'b010011111101: dataA <= 32'b00000101101101011111011101101010;
12'b010011111110: dataA <= 32'b01100111000011100110001100010110;
12'b010011111111: dataA <= 32'b00001110001000110100110110010000;
12'b010100000000: dataA <= 32'b10000010110101000100010100011000;
12'b010100000001: dataA <= 32'b00000101011101000110100000101100;
12'b010100000010: dataA <= 32'b00001011100101011101000010101010;
12'b010100000011: dataA <= 32'b00001010000100101111011101000101;
12'b010100000100: dataA <= 32'b10100100111111110100101101101111;
12'b010100000101: dataA <= 32'b00000110100110011010110010001010;
12'b010100000110: dataA <= 32'b10101111000111010100111010100101;
12'b010100000111: dataA <= 32'b00000001101010001010111111010110;
12'b010100001000: dataA <= 32'b00000000000010011110101000010110;
12'b010100001001: dataA <= 32'b00000000000000000000000000000000;
12'b010100001010: dataA <= 32'b01100111110011100110001011111100;
12'b010100001011: dataA <= 32'b00001000001001100011011010000000;
12'b010100001100: dataA <= 32'b01001001100111010001011100101011;
12'b010100001101: dataA <= 32'b00000011100011001000101001000110;
12'b010100001110: dataA <= 32'b11111101010001000010110011110000;
12'b010100001111: dataA <= 32'b00000110000001011000101011110011;
12'b010100010000: dataA <= 32'b01100111011011010100101010110010;
12'b010100010001: dataA <= 32'b00000101010010010001011110100000;
12'b010100010010: dataA <= 32'b01010001110101100010010101101110;
12'b010100010011: dataA <= 32'b00001011010110101101110101000001;
12'b010100010100: dataA <= 32'b11100101000010010000011001101000;
12'b010100010101: dataA <= 32'b00000110101001011011111010011010;
12'b010100010110: dataA <= 32'b01011011001000111011100001110011;
12'b010100010111: dataA <= 32'b00000110011001010010011101101011;
12'b010100011000: dataA <= 32'b01110010100000101100010001110111;
12'b010100011001: dataA <= 32'b00000100100010010101001111110011;
12'b010100011010: dataA <= 32'b01101000100010110001111001001100;
12'b010100011011: dataA <= 32'b00001001011110011100100111010101;
12'b010100011100: dataA <= 32'b01000100111000100001100001111000;
12'b010100011101: dataA <= 32'b00000101101001010000001100100010;
12'b010100011110: dataA <= 32'b11100111100101000010110000101100;
12'b010100011111: dataA <= 32'b00000101101011010011011111001110;
12'b010100100000: dataA <= 32'b01101011001010000100000111001010;
12'b010100100001: dataA <= 32'b00000101000001011011110110100011;
12'b010100100010: dataA <= 32'b11010101110111001001001010000001;
12'b010100100011: dataA <= 32'b00000110001100010110011101001010;
12'b010100100100: dataA <= 32'b00101111011101110101100110001001;
12'b010100100101: dataA <= 32'b00000100011100000111100011110101;
12'b010100100110: dataA <= 32'b01101100111010000001101000011101;
12'b010100100111: dataA <= 32'b00001000100001100011000011000101;
12'b010100101000: dataA <= 32'b11111101001110111000101011001000;
12'b010100101001: dataA <= 32'b00001010100100101010110011100001;
12'b010100101010: dataA <= 32'b00110001110011100110001000101001;
12'b010100101011: dataA <= 32'b00000100000111001110110011001011;
12'b010100101100: dataA <= 32'b10101010110010011100011000101100;
12'b010100101101: dataA <= 32'b00001100010111100111001011010011;
12'b010100101110: dataA <= 32'b00001010110001011000010101111000;
12'b010100101111: dataA <= 32'b00001111010100110001000000111100;
12'b010100110000: dataA <= 32'b10010111100001100000010111010000;
12'b010100110001: dataA <= 32'b00001011100010101111010101010011;
12'b010100110010: dataA <= 32'b01100011011100111100000100011011;
12'b010100110011: dataA <= 32'b00001100001110101111001110001100;
12'b010100110100: dataA <= 32'b11101000101010100000011001001000;
12'b010100110101: dataA <= 32'b00001000100111100001001111001001;
12'b010100110110: dataA <= 32'b11100100101010111110001001100100;
12'b010100110111: dataA <= 32'b00000011100111000111010110110101;
12'b010100111000: dataA <= 32'b10000100101101001000100100001010;
12'b010100111001: dataA <= 32'b00001001000101100011100101011100;
12'b010100111010: dataA <= 32'b00100110111010000101010111111101;
12'b010100111011: dataA <= 32'b00000110110101010111101011000011;
12'b010100111100: dataA <= 32'b01101100111000111101010001001000;
12'b010100111101: dataA <= 32'b00001011001001101111011110111010;
12'b010100111110: dataA <= 32'b11110101001110010001101000101011;
12'b010100111111: dataA <= 32'b00000100101001010101010111110010;
12'b010101000000: dataA <= 32'b01001011000101001110010010111010;
12'b010101000001: dataA <= 32'b00001101000110101011001000110101;
12'b010101000010: dataA <= 32'b01011000011100100001100011010010;
12'b010101000011: dataA <= 32'b00001001001101100101001001111111;
12'b010101000100: dataA <= 32'b00101101001001011001110101111011;
12'b010101000101: dataA <= 32'b00000101001011000110011110100001;
12'b010101000110: dataA <= 32'b01010000111101101100100110011000;
12'b010101000111: dataA <= 32'b00000100111101001111110001001010;
12'b010101001000: dataA <= 32'b00100000101000111001100001001010;
12'b010101001001: dataA <= 32'b00001101011010100000111110110111;
12'b010101001010: dataA <= 32'b01011111101001001011100011110011;
12'b010101001011: dataA <= 32'b00000100111010000101000001111000;
12'b010101001100: dataA <= 32'b01001101100001011101110011111010;
12'b010101001101: dataA <= 32'b00001011101010101001010101001111;
12'b010101001110: dataA <= 32'b01001100011110101100001010111100;
12'b010101001111: dataA <= 32'b00001001111000011110110101011011;
12'b010101010000: dataA <= 32'b01010101110111001001001100111011;
12'b010101010001: dataA <= 32'b00001001001000100010110101010101;
12'b010101010010: dataA <= 32'b11100001110101100001110110111001;
12'b010101010011: dataA <= 32'b00000110001100011011011101110010;
12'b010101010100: dataA <= 32'b01100111000011010110101011011000;
12'b010101010101: dataA <= 32'b00001111001010110110111110100000;
12'b010101010110: dataA <= 32'b00000100101000111011110011010110;
12'b010101010111: dataA <= 32'b00000011111100001010010100100100;
12'b010101011000: dataA <= 32'b10000111011101010100110011001000;
12'b010101011001: dataA <= 32'b00001011000101101011100001000100;
12'b010101011010: dataA <= 32'b10100100111111101101011101110001;
12'b010101011011: dataA <= 32'b00000111100110011100110010010010;
12'b010101011100: dataA <= 32'b00101111001111001101011011100110;
12'b010101011101: dataA <= 32'b00000010101000001010110011000111;
12'b010101011110: dataA <= 32'b00000000000010001110100111110110;
12'b010101011111: dataA <= 32'b00000000000000000000000000000000;
12'b010101100000: dataA <= 32'b11111000110011000000111110001000;
12'b010101100001: dataA <= 32'b00000100101111101100111000001011;
12'b010101100010: dataA <= 32'b11110011101100101001010101100110;
12'b010101100011: dataA <= 32'b00000001111000010101101111001101;
12'b010101100100: dataA <= 32'b01101000000101011101111000011000;
12'b010101100101: dataA <= 32'b00000000110011010101001101111000;
12'b010101100110: dataA <= 32'b11101100110010010001011001001010;
12'b010101100111: dataA <= 32'b00001001010101101111011100001010;
12'b010101101000: dataA <= 32'b11111011011101001100110111010100;
12'b010101101001: dataA <= 32'b00001011001001111010100100101101;
12'b010101101010: dataA <= 32'b00100000110100001011010100001100;
12'b010101101011: dataA <= 32'b00000100110010111101001001011011;
12'b010101101100: dataA <= 32'b10100101001001110110001001111100;
12'b010101101101: dataA <= 32'b00001100110011001111011001101100;
12'b010101101110: dataA <= 32'b01010000011010001110101011111100;
12'b010101101111: dataA <= 32'b00000001010110100111010101101000;
12'b010101110000: dataA <= 32'b01010000101100111010010110001101;
12'b010101110001: dataA <= 32'b00001111001101010011000110101001;
12'b010101110010: dataA <= 32'b11011101110100110110111100011100;
12'b010101110011: dataA <= 32'b00000100110100000111011101001110;
12'b010101110100: dataA <= 32'b10110010110001011101110110011110;
12'b010101110101: dataA <= 32'b00000101110100101111011011011001;
12'b010101110110: dataA <= 32'b11100100101010000011110101010001;
12'b010101110111: dataA <= 32'b00000000110101111011001001101010;
12'b010101111000: dataA <= 32'b10111011010100100001100000101011;
12'b010101111001: dataA <= 32'b00000110010011001111010001011101;
12'b010101111010: dataA <= 32'b01101110100010110100010100110011;
12'b010101111011: dataA <= 32'b00001110010111110001110010100000;
12'b010101111100: dataA <= 32'b11011100100100110011111110101111;
12'b010101111101: dataA <= 32'b00000000101110100000111010101001;
12'b010101111110: dataA <= 32'b11100110000100010010000100001001;
12'b010101111111: dataA <= 32'b00000010001010011000101000111000;
12'b010110000000: dataA <= 32'b10111000011111000000110100101110;
12'b010110000001: dataA <= 32'b00000011110111011001100001100001;
12'b010110000010: dataA <= 32'b01011000101010001011000110001110;
12'b010110000011: dataA <= 32'b00001011100111100100110001110001;
12'b010110000100: dataA <= 32'b00011001101000001101001100010100;
12'b010110000101: dataA <= 32'b00001010000001100000011110000110;
12'b010110000110: dataA <= 32'b01110001010000001100111000010001;
12'b010110000111: dataA <= 32'b00000001001000101010100001110101;
12'b010110001000: dataA <= 32'b10101110111010000110001101110111;
12'b010110001001: dataA <= 32'b00000111000111100110100010001011;
12'b010110001010: dataA <= 32'b10010100101100001010110100001101;
12'b010110001011: dataA <= 32'b00000011101110100110111100111001;
12'b010110001100: dataA <= 32'b01010100110111000010000010001100;
12'b010110001101: dataA <= 32'b00000011111000101011110010111010;
12'b010110001110: dataA <= 32'b00010111110100010101100101010111;
12'b010110001111: dataA <= 32'b00000010101101110010111010010101;
12'b010110010000: dataA <= 32'b11011100110010101011111110110000;
12'b010110010001: dataA <= 32'b00001010110010110101010001100001;
12'b010110010010: dataA <= 32'b00011100100110101110000100011101;
12'b010110010011: dataA <= 32'b00000100101001101110100001001010;
12'b010110010100: dataA <= 32'b01100110010100110011010101101110;
12'b010110010101: dataA <= 32'b00000100110110101011010101011000;
12'b010110010110: dataA <= 32'b01100011101011001101101101011010;
12'b010110010111: dataA <= 32'b00000011000101100100101010101110;
12'b010110011000: dataA <= 32'b00001111001100110110111001011001;
12'b010110011001: dataA <= 32'b00000110101101100100110111101100;
12'b010110011010: dataA <= 32'b11100100100100111101001101110100;
12'b010110011011: dataA <= 32'b00000101110101001111110000100010;
12'b010110011100: dataA <= 32'b10011111011110010100101100010011;
12'b010110011101: dataA <= 32'b00001110110110111001100001001101;
12'b010110011110: dataA <= 32'b01010100111100110110000101011101;
12'b010110011111: dataA <= 32'b00001101000101011110111111100010;
12'b010110100000: dataA <= 32'b00110101000001110101101001111000;
12'b010110100001: dataA <= 32'b00001101010110100001110100001100;
12'b010110100010: dataA <= 32'b10110001100110111101001101011000;
12'b010110100011: dataA <= 32'b00000101001000101010101111101101;
12'b010110100100: dataA <= 32'b00001111100110000010101110001010;
12'b010110100101: dataA <= 32'b00001100001100011011000001101101;
12'b010110100110: dataA <= 32'b01111011010100100001101101100110;
12'b010110100111: dataA <= 32'b00000100001101011010111010101101;
12'b010110101000: dataA <= 32'b01111010111100111100111100110010;
12'b010110101001: dataA <= 32'b00000110010011101111001001011100;
12'b010110101010: dataA <= 32'b11100000110011010001011100001001;
12'b010110101011: dataA <= 32'b00000101000001011110010000001010;
12'b010110101100: dataA <= 32'b11010101110101111110001011011001;
12'b010110101101: dataA <= 32'b00001110011000001011101010000110;
12'b010110101110: dataA <= 32'b11101111110010011101010100011001;
12'b010110101111: dataA <= 32'b00000010101001110000101010010101;
12'b010110110000: dataA <= 32'b01011110110110101000101000100100;
12'b010110110001: dataA <= 32'b00000011010000011001000101010011;
12'b010110110010: dataA <= 32'b11100110100010101001100011001000;
12'b010110110011: dataA <= 32'b00000100011010011001101011100001;
12'b010110110100: dataA <= 32'b00000000000011010011101011010000;
12'b010110110101: dataA <= 32'b00000000000000000000000000000000;
12'b010110110110: dataA <= 32'b10110110101010110000101101100101;
12'b010110110111: dataA <= 32'b00000100110000101100110100001100;
12'b010110111000: dataA <= 32'b01110111100100100010000100100111;
12'b010110111001: dataA <= 32'b00000010111011011001110011010101;
12'b010110111010: dataA <= 32'b01100010000101101110001001011000;
12'b010110111011: dataA <= 32'b00000001010110010111010001100000;
12'b010110111100: dataA <= 32'b10101010101101111001011000101010;
12'b010110111101: dataA <= 32'b00001001110101110011010100001011;
12'b010110111110: dataA <= 32'b00111101010001010101000111110100;
12'b010110111111: dataA <= 32'b00001010001000111000011100111110;
12'b010111000000: dataA <= 32'b01100000110100001100000100001110;
12'b010111000001: dataA <= 32'b00000100110011111100111101011011;
12'b010111000010: dataA <= 32'b10100101001010000110001010111011;
12'b010111000011: dataA <= 32'b00001100110001010011100001101100;
12'b010111000100: dataA <= 32'b01001100100010011110101100111010;
12'b010111000101: dataA <= 32'b00000010011001101001010001010000;
12'b010111000110: dataA <= 32'b00001110110100110010110110001110;
12'b010111000111: dataA <= 32'b00001111001010010011001010011001;
12'b010111001000: dataA <= 32'b00100001110101000111011101011010;
12'b010111001001: dataA <= 32'b00000101010101001001101001011111;
12'b010111001010: dataA <= 32'b00110000101001101110000111111110;
12'b010111001011: dataA <= 32'b00000110010101110001010011001001;
12'b010111001100: dataA <= 32'b11100010101010000011110101010010;
12'b010111001101: dataA <= 32'b00000001110111111011000001100010;
12'b010111001110: dataA <= 32'b11111101001000010010000000101101;
12'b010111001111: dataA <= 32'b00000110110100010001011001100101;
12'b010111010000: dataA <= 32'b01101010011010110100000101010100;
12'b010111010001: dataA <= 32'b00001111010100110101101010010000;
12'b010111010010: dataA <= 32'b10011010100100111100011110001101;
12'b010111010011: dataA <= 32'b00000000110001100000111010011001;
12'b010111010100: dataA <= 32'b01100000000100001010110011101011;
12'b010111010101: dataA <= 32'b00000001101100010110101100100001;
12'b010111010110: dataA <= 32'b11110100010010110000100100101111;
12'b010111010111: dataA <= 32'b00000100111001011101100001010001;
12'b010111011000: dataA <= 32'b01010110101110001011000110001110;
12'b010111011001: dataA <= 32'b00001010100110100010110001100001;
12'b010111011010: dataA <= 32'b00011101101100010101111100110010;
12'b010111011011: dataA <= 32'b00001000100001011100100010010110;
12'b010111011100: dataA <= 32'b01110011001000010101101000010001;
12'b010111011101: dataA <= 32'b00000000101011100110011101111101;
12'b010111011110: dataA <= 32'b10101110110010010110001110110101;
12'b010111011111: dataA <= 32'b00000110000111100010100010001011;
12'b010111100000: dataA <= 32'b00010010110000001011010100001111;
12'b010111100001: dataA <= 32'b00000011110000100110111000101010;
12'b010111100010: dataA <= 32'b11010100111010110001100010001110;
12'b010111100011: dataA <= 32'b00000100111010101111101110101001;
12'b010111100100: dataA <= 32'b00011101111000100110010110011000;
12'b010111100101: dataA <= 32'b00000010110000110010110010011101;
12'b010111100110: dataA <= 32'b00011010110010101011101110101110;
12'b010111100111: dataA <= 32'b00001010110001110111001001010010;
12'b010111101000: dataA <= 32'b10011010100110111101110101111110;
12'b010111101001: dataA <= 32'b00000100001011101010011000111010;
12'b010111101010: dataA <= 32'b10100010010000110011110101101111;
12'b010111101011: dataA <= 32'b00000101110111101101010001000000;
12'b010111101100: dataA <= 32'b00100111101011010101001110010111;
12'b010111101101: dataA <= 32'b00000010100111100010101010111110;
12'b010111101110: dataA <= 32'b10010001010101000111001010011000;
12'b010111101111: dataA <= 32'b00000110101101100100110111101011;
12'b010111110000: dataA <= 32'b01100010100101000101101110010010;
12'b010111110001: dataA <= 32'b00000110010110010101110100011011;
12'b010111110010: dataA <= 32'b11100011011010010100101100010001;
12'b010111110011: dataA <= 32'b00001111010011111011011001011101;
12'b010111110100: dataA <= 32'b11010101000001000110100110111110;
12'b010111110101: dataA <= 32'b00001100000011011110111111010001;
12'b010111110110: dataA <= 32'b11110010111001111101101010110111;
12'b010111110111: dataA <= 32'b00001101110100100101110000001100;
12'b010111111000: dataA <= 32'b11110101011111000100101110010110;
12'b010111111001: dataA <= 32'b00000100001001101000101011110100;
12'b010111111010: dataA <= 32'b00010101101101111010101101101000;
12'b010111111011: dataA <= 32'b00001011101010011011000001110101;
12'b010111111100: dataA <= 32'b00111101001000010010001100100100;
12'b010111111101: dataA <= 32'b00000100001111011010111010110101;
12'b010111111110: dataA <= 32'b10111000110101000101011100110000;
12'b010111111111: dataA <= 32'b00000110110100101111000001011100;
12'b011000000000: dataA <= 32'b01100000110011000000111011000111;
12'b011000000001: dataA <= 32'b00000100000011011010010100001011;
12'b011000000010: dataA <= 32'b10011011111010001101111100010111;
12'b011000000011: dataA <= 32'b00001110110101010001110010010110;
12'b011000000100: dataA <= 32'b11110011101010100101000101011010;
12'b011000000101: dataA <= 32'b00000010001011101110100010100101;
12'b011000000110: dataA <= 32'b10011110110110010000010111100100;
12'b011000000111: dataA <= 32'b00000011010010011001001001010011;
12'b011000001000: dataA <= 32'b01100010100010011001010010101010;
12'b011000001001: dataA <= 32'b00000101011100011111101011010001;
12'b011000001010: dataA <= 32'b00000000000011010011001011001111;
12'b011000001011: dataA <= 32'b00000000000000000000000000000000;
12'b011000001100: dataA <= 32'b01110100100010011000011100000011;
12'b011000001101: dataA <= 32'b00000101010001101010101100001101;
12'b011000001110: dataA <= 32'b10111001011100010010100011101001;
12'b011000001111: dataA <= 32'b00000100011100011111110111011100;
12'b011000010000: dataA <= 32'b10011100000101110110001010010111;
12'b011000010001: dataA <= 32'b00000001111000011001010101001000;
12'b011000010010: dataA <= 32'b01101000101001101001011000001010;
12'b011000010011: dataA <= 32'b00001010010100110011001100001100;
12'b011000010100: dataA <= 32'b10111101000101011101011000010100;
12'b011000010101: dataA <= 32'b00001001100111110100010101001110;
12'b011000010110: dataA <= 32'b10011110110100001100110011101111;
12'b011000010111: dataA <= 32'b00000101010101111100110001010011;
12'b011000011000: dataA <= 32'b11100111000110010101111011111010;
12'b011000011001: dataA <= 32'b00001100101111010101100101110100;
12'b011000011010: dataA <= 32'b11001010101010101110011101111000;
12'b011000011011: dataA <= 32'b00000011011011101011001101000000;
12'b011000011100: dataA <= 32'b11001110111000101011010101101110;
12'b011000011101: dataA <= 32'b00001110001000010101010010001000;
12'b011000011110: dataA <= 32'b01100111110001011111101110011000;
12'b011000011111: dataA <= 32'b00000101110110001111110001110111;
12'b011000100000: dataA <= 32'b11101110100001110110001001011110;
12'b011000100001: dataA <= 32'b00000110110101110011001010111000;
12'b011000100010: dataA <= 32'b00100000101010000011110101110011;
12'b011000100011: dataA <= 32'b00000010111010111010110101011011;
12'b011000100100: dataA <= 32'b11111101000000001010110000110000;
12'b011000100101: dataA <= 32'b00000110110100010011011101110101;
12'b011000100110: dataA <= 32'b01100110011010110011100101110101;
12'b011000100111: dataA <= 32'b00001111010010111001100001111000;
12'b011000101000: dataA <= 32'b10010110101000111100111101101010;
12'b011000101001: dataA <= 32'b00000000110100100000111010001001;
12'b011000101010: dataA <= 32'b00011010000100001011100011001101;
12'b011000101011: dataA <= 32'b00000001001111010100110000011010;
12'b011000101100: dataA <= 32'b00101110001110011000010100110001;
12'b011000101101: dataA <= 32'b00000101111010100001100001000010;
12'b011000101110: dataA <= 32'b10010100110010000011000110001111;
12'b011000101111: dataA <= 32'b00001001100101100010101101010001;
12'b011000110000: dataA <= 32'b11100001101100100110011100110000;
12'b011000110001: dataA <= 32'b00000111000001011010100010100101;
12'b011000110010: dataA <= 32'b01110011000000011110001000010001;
12'b011000110011: dataA <= 32'b00000000101110100010011010000101;
12'b011000110100: dataA <= 32'b10101100101110100101111110110010;
12'b011000110101: dataA <= 32'b00000101001000100000011110001011;
12'b011000110110: dataA <= 32'b10010010110100001100000100010000;
12'b011000110111: dataA <= 32'b00000100010010100110111000100010;
12'b011000111000: dataA <= 32'b10010100111110100001010001110000;
12'b011000111001: dataA <= 32'b00000101111011110011100110100001;
12'b011000111010: dataA <= 32'b11100001111000110110110111011001;
12'b011000111011: dataA <= 32'b00000010110010110000101010100100;
12'b011000111100: dataA <= 32'b01011010110010101011011110001011;
12'b011000111101: dataA <= 32'b00001010110000110111000001001010;
12'b011000111110: dataA <= 32'b11010110101011000101010111011110;
12'b011000111111: dataA <= 32'b00000011101100100110011000110010;
12'b011001000000: dataA <= 32'b00011110010000110100010101110000;
12'b011001000001: dataA <= 32'b00000110011000101111001000110001;
12'b011001000010: dataA <= 32'b10101011100111011100011111010101;
12'b011001000011: dataA <= 32'b00000001101010100000101011001101;
12'b011001000100: dataA <= 32'b11010011011001011111101011010111;
12'b011001000101: dataA <= 32'b00000110001110100010110011100010;
12'b011001000110: dataA <= 32'b11011110100101001101111110010000;
12'b011001000111: dataA <= 32'b00000110110110011001111000011011;
12'b011001001000: dataA <= 32'b00100101011010011100011100001111;
12'b011001001001: dataA <= 32'b00001111010000111101001101100110;
12'b011001001010: dataA <= 32'b01010111000101010110110111111110;
12'b011001001011: dataA <= 32'b00001011000010011110111111001001;
12'b011001001100: dataA <= 32'b10110010110010001101101011010110;
12'b011001001101: dataA <= 32'b00001110010010101011101100010101;
12'b011001001110: dataA <= 32'b00110111010111000100011110110100;
12'b011001001111: dataA <= 32'b00000011101011100110100111110100;
12'b011001010000: dataA <= 32'b00011001110001110010111100100110;
12'b011001010001: dataA <= 32'b00001011001001011011000101111101;
12'b011001010010: dataA <= 32'b10111100111100001010111011100011;
12'b011001010011: dataA <= 32'b00000100010000011010111110111100;
12'b011001010100: dataA <= 32'b11110110101001001101101100101110;
12'b011001010101: dataA <= 32'b00000110110100101110111101100100;
12'b011001010110: dataA <= 32'b00011110110010101000101010100110;
12'b011001010111: dataA <= 32'b00000010100101010110010100001100;
12'b011001011000: dataA <= 32'b10011111111010010101111101010101;
12'b011001011001: dataA <= 32'b00001111010011010101111010100110;
12'b011001011010: dataA <= 32'b10110111100010101100110110111011;
12'b011001011011: dataA <= 32'b00000001101101101010011110101101;
12'b011001011100: dataA <= 32'b11011100110101111000010110100100;
12'b011001011101: dataA <= 32'b00000011110100011001001001010011;
12'b011001011110: dataA <= 32'b11100000011110001001010010001101;
12'b011001011111: dataA <= 32'b00000110011101100011101011000000;
12'b011001100000: dataA <= 32'b00000000000011001010101010101110;
12'b011001100001: dataA <= 32'b00000000000000000000000000000000;
12'b011001100010: dataA <= 32'b11110000011010000000011011000010;
12'b011001100011: dataA <= 32'b00000101010011101000101000011101;
12'b011001100100: dataA <= 32'b00111101010000010011010011001010;
12'b011001100101: dataA <= 32'b00000101011110100011110011100100;
12'b011001100110: dataA <= 32'b11010110000110000110001010110110;
12'b011001100111: dataA <= 32'b00000010111010011011011000111000;
12'b011001101000: dataA <= 32'b00100110100101011001100111101010;
12'b011001101001: dataA <= 32'b00001010110011110101000100001101;
12'b011001101010: dataA <= 32'b11111100111001100101101000010100;
12'b011001101011: dataA <= 32'b00001000100110101110001101011110;
12'b011001101100: dataA <= 32'b11011110110100010101100100010001;
12'b011001101101: dataA <= 32'b00000101110101111010100101010011;
12'b011001101110: dataA <= 32'b11100111000110011101111100111000;
12'b011001101111: dataA <= 32'b00001100101101011001101001110100;
12'b011001110000: dataA <= 32'b01001000110010110110001110010110;
12'b011001110001: dataA <= 32'b00000100011101101101001000101001;
12'b011001110010: dataA <= 32'b11001111000000101011110101101111;
12'b011001110011: dataA <= 32'b00001101000101010111010101111000;
12'b011001110100: dataA <= 32'b01101011101101110111101110110101;
12'b011001110101: dataA <= 32'b00000110110111010011110110000111;
12'b011001110110: dataA <= 32'b01101010011110000110001010111110;
12'b011001110111: dataA <= 32'b00000111010110110011000010100000;
12'b011001111000: dataA <= 32'b01011110101010000011110101110100;
12'b011001111001: dataA <= 32'b00000011111100111000101001011011;
12'b011001111010: dataA <= 32'b11111100110100001011100000110011;
12'b011001111011: dataA <= 32'b00000111010100010111100001111101;
12'b011001111100: dataA <= 32'b01100010010110101011010110010110;
12'b011001111101: dataA <= 32'b00001111001111111011010101100000;
12'b011001111110: dataA <= 32'b10010100101101000101001101001000;
12'b011001111111: dataA <= 32'b00000001010111100000111001111001;
12'b011010000000: dataA <= 32'b10010100000100001100010011001111;
12'b011010000001: dataA <= 32'b00000001110001010010110100001010;
12'b011010000010: dataA <= 32'b10101010000110000000010101010010;
12'b011010000011: dataA <= 32'b00000110111011100011100000111010;
12'b011010000100: dataA <= 32'b11010010110101111011000110010000;
12'b011010000101: dataA <= 32'b00001000100100100000101101001001;
12'b011010000110: dataA <= 32'b10100101101000110110111100101110;
12'b011010000111: dataA <= 32'b00000101100001010110100110101101;
12'b011010001000: dataA <= 32'b01110010111000101110101000110001;
12'b011010001001: dataA <= 32'b00000000110001100000011010001101;
12'b011010001010: dataA <= 32'b01101010101010101101101111001111;
12'b011010001011: dataA <= 32'b00000100101001011100100010000011;
12'b011010001100: dataA <= 32'b01010000111100001100110100010010;
12'b011010001101: dataA <= 32'b00000100010011100110110100011011;
12'b011010001110: dataA <= 32'b10010101000010010001000010010011;
12'b011010001111: dataA <= 32'b00000111011011110111011110010001;
12'b011010010000: dataA <= 32'b10100111110101000111010111111001;
12'b011010010001: dataA <= 32'b00000011010100101110100010100100;
12'b011010010010: dataA <= 32'b10011000110110100011001101101001;
12'b011010010011: dataA <= 32'b00001010101111110110111000111010;
12'b011010010100: dataA <= 32'b01010100101111001100111000111110;
12'b011010010101: dataA <= 32'b00000011001110100010010100110011;
12'b011010010110: dataA <= 32'b10011010010100111100110101110000;
12'b011010010111: dataA <= 32'b00000111011001101111000100100001;
12'b011010011000: dataA <= 32'b00101101100011011011111111010010;
12'b011010011001: dataA <= 32'b00000001001100011110101011010101;
12'b011010011010: dataA <= 32'b01010101100001101111101011110110;
12'b011010011011: dataA <= 32'b00000110001110100010110011011010;
12'b011010011100: dataA <= 32'b10011100100101011110001110001101;
12'b011010011101: dataA <= 32'b00000111110111011111111000011100;
12'b011010011110: dataA <= 32'b01100111011010011100011100001110;
12'b011010011111: dataA <= 32'b00001111001101111101000001110110;
12'b011010100000: dataA <= 32'b11010111001001101111001001011110;
12'b011010100001: dataA <= 32'b00001001100001011110111110110000;
12'b011010100010: dataA <= 32'b00110000101010010101011100010101;
12'b011010100011: dataA <= 32'b00001110001111101111101000011110;
12'b011010100100: dataA <= 32'b01111001001011000011111111010001;
12'b011010100101: dataA <= 32'b00000011101100100100100111110011;
12'b011010100110: dataA <= 32'b00011101110001101010111011100100;
12'b011010100111: dataA <= 32'b00001010100111011011000110000101;
12'b011010101000: dataA <= 32'b01111100110100001011101010000001;
12'b011010101001: dataA <= 32'b00000100010010011010111110111100;
12'b011010101010: dataA <= 32'b11110100100001010110001100001100;
12'b011010101011: dataA <= 32'b00000111010100101110110101100100;
12'b011010101100: dataA <= 32'b11011100110110010000011001100101;
12'b011010101101: dataA <= 32'b00000001100111010010011000001100;
12'b011010101110: dataA <= 32'b01100101111010100101101101010011;
12'b011010101111: dataA <= 32'b00001111010000011011111010110110;
12'b011010110000: dataA <= 32'b00111001011010110100100111111100;
12'b011010110001: dataA <= 32'b00000001110000100110011010110101;
12'b011010110010: dataA <= 32'b00011100110101101000010101100101;
12'b011010110011: dataA <= 32'b00000100010110011011001101010100;
12'b011010110100: dataA <= 32'b10011100100001110001010001101111;
12'b011010110101: dataA <= 32'b00000111111101100111101010101000;
12'b011010110110: dataA <= 32'b00000000000011000010011010101100;
12'b011010110111: dataA <= 32'b00000000000000000000000000000000;
12'b011010111000: dataA <= 32'b10101100010001101000011001100001;
12'b011010111001: dataA <= 32'b00000101110100100110100100101110;
12'b011010111010: dataA <= 32'b10111101001000001011110010101100;
12'b011010111011: dataA <= 32'b00000110111110101001110011011011;
12'b011010111100: dataA <= 32'b01010000001010010110001011010101;
12'b011010111101: dataA <= 32'b00000100011100011101011000101001;
12'b011010111110: dataA <= 32'b11100100100001010001110111001010;
12'b011010111111: dataA <= 32'b00001010110010110100111100010101;
12'b011011000000: dataA <= 32'b00111100101101101101111000110100;
12'b011011000001: dataA <= 32'b00000111100110101010000101101111;
12'b011011000010: dataA <= 32'b00011110110100011110000100010010;
12'b011011000011: dataA <= 32'b00000110110110111000011101010100;
12'b011011000100: dataA <= 32'b11100111000010100101101101110110;
12'b011011000101: dataA <= 32'b00001100001011011101101001111100;
12'b011011000110: dataA <= 32'b11000110111111000101101110110011;
12'b011011000111: dataA <= 32'b00000101111110101101000100011001;
12'b011011001000: dataA <= 32'b00001111001000101100010101110000;
12'b011011001001: dataA <= 32'b00001100000011011001011001100001;
12'b011011001010: dataA <= 32'b01110001101010001111101111010010;
12'b011011001011: dataA <= 32'b00000111010111011001111010011111;
12'b011011001100: dataA <= 32'b01101000011010010110001011111100;
12'b011011001101: dataA <= 32'b00000111110110110010111110010000;
12'b011011001110: dataA <= 32'b10011100101010000011110110010101;
12'b011011001111: dataA <= 32'b00000100111101110110100001010011;
12'b011011010000: dataA <= 32'b11111010101000001100010001010110;
12'b011011010001: dataA <= 32'b00000111110100011011100110001101;
12'b011011010010: dataA <= 32'b10011110010110101011000110110111;
12'b011011010011: dataA <= 32'b00001111001100111101001001001000;
12'b011011010100: dataA <= 32'b10010010110001001101101100100110;
12'b011011010101: dataA <= 32'b00000010011001011110111001101001;
12'b011011010110: dataA <= 32'b01010000001100001101000011010000;
12'b011011010111: dataA <= 32'b00000001110100010010111000001011;
12'b011011011000: dataA <= 32'b11100100000101101000010101010011;
12'b011011011001: dataA <= 32'b00000111111011100111100000110010;
12'b011011011010: dataA <= 32'b01010010111001110011000110010001;
12'b011011011011: dataA <= 32'b00000111000100011110101100111010;
12'b011011011100: dataA <= 32'b01101001101001000111011100001100;
12'b011011011101: dataA <= 32'b00000100000010010100101010110101;
12'b011011011110: dataA <= 32'b00110000110001000111001000110001;
12'b011011011111: dataA <= 32'b00000000110100011100011010010101;
12'b011011100000: dataA <= 32'b01101000100110110101011110101101;
12'b011011100001: dataA <= 32'b00000100001011011010100010000011;
12'b011011100010: dataA <= 32'b11010001000000010101100100110011;
12'b011011100011: dataA <= 32'b00000100110100100100110000011011;
12'b011011100100: dataA <= 32'b10010101000110000001000010110101;
12'b011011100101: dataA <= 32'b00001000011100111001010110000001;
12'b011011100110: dataA <= 32'b01101101110001011111101000111001;
12'b011011100111: dataA <= 32'b00000011110101101010011110101100;
12'b011011101000: dataA <= 32'b00011000111010011010111100100111;
12'b011011101001: dataA <= 32'b00001010101110110100110000111011;
12'b011011101010: dataA <= 32'b11010010110011010100011010011110;
12'b011011101011: dataA <= 32'b00000011010000011110010100110011;
12'b011011101100: dataA <= 32'b00010110010100111101010101110001;
12'b011011101101: dataA <= 32'b00001000011001101110111100010010;
12'b011011101110: dataA <= 32'b10110001011011011011011111001111;
12'b011011101111: dataA <= 32'b00000001001111011100101011010100;
12'b011011110000: dataA <= 32'b11011001100010000111101100010100;
12'b011011110001: dataA <= 32'b00000110001111100000110011001001;
12'b011011110010: dataA <= 32'b00011010100101101110011101101011;
12'b011011110011: dataA <= 32'b00001000010111100101111000100101;
12'b011011110100: dataA <= 32'b01101001010110011100001100001100;
12'b011011110101: dataA <= 32'b00001111001011111100110110000110;
12'b011011110110: dataA <= 32'b10011001001101111111001010111101;
12'b011011110111: dataA <= 32'b00001000000001011110111110100000;
12'b011011111000: dataA <= 32'b10101110100010011101011100010011;
12'b011011111001: dataA <= 32'b00001110001101110011100100101110;
12'b011011111010: dataA <= 32'b11111001000011000011011111001110;
12'b011011111011: dataA <= 32'b00000011001110100000100011110010;
12'b011011111100: dataA <= 32'b00100011110001100011001010100011;
12'b011011111101: dataA <= 32'b00001001100111011101001010001101;
12'b011011111110: dataA <= 32'b11111010101000001100011001000001;
12'b011011111111: dataA <= 32'b00000100110011011011000010111011;
12'b011100000000: dataA <= 32'b00110010011001100110001100001010;
12'b011100000001: dataA <= 32'b00000111110100101100110001101101;
12'b011100000010: dataA <= 32'b10011100110101111000011000100101;
12'b011100000011: dataA <= 32'b00000001001001010000100000010101;
12'b011100000100: dataA <= 32'b11101011110110101101011101110001;
12'b011100000101: dataA <= 32'b00001111001101100001111010111101;
12'b011100000110: dataA <= 32'b11111011001110110100011000111011;
12'b011100000111: dataA <= 32'b00000001110010100010010110111100;
12'b011100001000: dataA <= 32'b01011010111001010000100100100110;
12'b011100001001: dataA <= 32'b00000100110111011101001101010100;
12'b011100001010: dataA <= 32'b01011010100001100001010010010001;
12'b011100001011: dataA <= 32'b00001001011101101011100110010000;
12'b011100001100: dataA <= 32'b00000000000010110001111010001011;
12'b011100001101: dataA <= 32'b00000000000000000000000000000000;
12'b011100001110: dataA <= 32'b00101000001101010000011000000001;
12'b011100001111: dataA <= 32'b00000110010100100100100100111111;
12'b011100010000: dataA <= 32'b11111100111100010100100010101110;
12'b011100010001: dataA <= 32'b00001000011110101101101111011010;
12'b011100010010: dataA <= 32'b00001100010010011101111011110100;
12'b011100010011: dataA <= 32'b00000101011110011111011000011010;
12'b011100010100: dataA <= 32'b01100000100001000010000110101010;
12'b011100010101: dataA <= 32'b00001011010001110100110100100110;
12'b011100010110: dataA <= 32'b00111010100001111101111001010011;
12'b011100010111: dataA <= 32'b00000111000110100100000110000111;
12'b011100011000: dataA <= 32'b01011100111000101110100100110100;
12'b011100011001: dataA <= 32'b00000111010111110100010101010100;
12'b011100011010: dataA <= 32'b11100110111110110101011110010100;
12'b011100011011: dataA <= 32'b00001011101001100011101010000100;
12'b011100011100: dataA <= 32'b01000111000111001101011111010000;
12'b011100011101: dataA <= 32'b00000111011110101101000000010010;
12'b011100011110: dataA <= 32'b01010001001100110100110101110001;
12'b011100011111: dataA <= 32'b00001011000010011011011001010001;
12'b011100100000: dataA <= 32'b00110101100010100111101111001111;
12'b011100100001: dataA <= 32'b00001000011000011111111010101111;
12'b011100100010: dataA <= 32'b01100100010110011101111101011010;
12'b011100100011: dataA <= 32'b00001000110110110010110101111000;
12'b011100100100: dataA <= 32'b11011010101010000011110111010101;
12'b011100100101: dataA <= 32'b00000110011110110010011001010011;
12'b011100100110: dataA <= 32'b11111000011100001101000001111000;
12'b011100100111: dataA <= 32'b00001000010100011111100110010101;
12'b011100101000: dataA <= 32'b11011010010110100010110111110111;
12'b011100101001: dataA <= 32'b00001110101001111100111100111000;
12'b011100101010: dataA <= 32'b10010010110101010101111011100101;
12'b011100101011: dataA <= 32'b00000011011011011110111001011001;
12'b011100101100: dataA <= 32'b00001010010100010101110011010010;
12'b011100101101: dataA <= 32'b00000010010110010010111100001100;
12'b011100101110: dataA <= 32'b01011110000101010000010101110100;
12'b011100101111: dataA <= 32'b00001000111011101011011100101011;
12'b011100110000: dataA <= 32'b10010010111101110011000110010001;
12'b011100110001: dataA <= 32'b00000110000101011100101100110010;
12'b011100110010: dataA <= 32'b00101101100101011111101100001011;
12'b011100110011: dataA <= 32'b00000011000100010010101110111101;
12'b011100110100: dataA <= 32'b00110000101101010111101000110000;
12'b011100110101: dataA <= 32'b00000001010111011000011110011101;
12'b011100110110: dataA <= 32'b01100100100010111101001110101010;
12'b011100110111: dataA <= 32'b00000011101100010110100110000011;
12'b011100111000: dataA <= 32'b10010011001000011110000101010100;
12'b011100111001: dataA <= 32'b00000101010110100010110000011100;
12'b011100111010: dataA <= 32'b10010101001001110001000011010111;
12'b011100111011: dataA <= 32'b00001001011011111011001001110001;
12'b011100111100: dataA <= 32'b00110001101101110111101001111000;
12'b011100111101: dataA <= 32'b00000100010111100110011010101100;
12'b011100111110: dataA <= 32'b10011000111010010010101011100101;
12'b011100111111: dataA <= 32'b00001010101101110100101000110011;
12'b011101000000: dataA <= 32'b01010010110111010011111011011101;
12'b011101000001: dataA <= 32'b00000011010001011010010100110100;
12'b011101000010: dataA <= 32'b11010010011001001101100110010010;
12'b011101000011: dataA <= 32'b00001000111001101110111000001010;
12'b011101000100: dataA <= 32'b00110011010111010010111111001100;
12'b011101000101: dataA <= 32'b00000001010001011010101011011100;
12'b011101000110: dataA <= 32'b01011101100110011111101100110010;
12'b011101000111: dataA <= 32'b00000110010000011110110010111001;
12'b011101001000: dataA <= 32'b10011000101001111110011101001001;
12'b011101001001: dataA <= 32'b00001001010110101011110100101101;
12'b011101001010: dataA <= 32'b01101011010010011011111011101010;
12'b011101001011: dataA <= 32'b00001110001000111100101010001110;
12'b011101001100: dataA <= 32'b10011001001110010111001100011100;
12'b011101001101: dataA <= 32'b00000110100001011110111110001000;
12'b011101001110: dataA <= 32'b00101010011110100101001100110001;
12'b011101001111: dataA <= 32'b00001101101010110101011101000111;
12'b011101010000: dataA <= 32'b00111000110110111011001110101011;
12'b011101010001: dataA <= 32'b00000011010000011110100011100010;
12'b011101010010: dataA <= 32'b00100111110001100011001001000010;
12'b011101010011: dataA <= 32'b00001000100110011101001010010101;
12'b011101010100: dataA <= 32'b10111000011100001101000111100001;
12'b011101010101: dataA <= 32'b00000101010100011011000010111011;
12'b011101010110: dataA <= 32'b00101110010101110110011011001001;
12'b011101010111: dataA <= 32'b00001000010100101010101101110101;
12'b011101011000: dataA <= 32'b00011010110101100000010111000101;
12'b011101011001: dataA <= 32'b00000000101100001100100100011110;
12'b011101011010: dataA <= 32'b10110001110010110101001101101111;
12'b011101011011: dataA <= 32'b00001110101010100111111011001101;
12'b011101011100: dataA <= 32'b10111101000010110100001010011011;
12'b011101011101: dataA <= 32'b00000010010101011110010110111100;
12'b011101011110: dataA <= 32'b10011010111000111000110011101000;
12'b011101011111: dataA <= 32'b00000101111000011101001101010100;
12'b011101100000: dataA <= 32'b01010110100101010001100010010100;
12'b011101100001: dataA <= 32'b00001010011100101101100010000000;
12'b011101100010: dataA <= 32'b00000000000010101001101001101011;
12'b011101100011: dataA <= 32'b00000000000000000000000000000000;
12'b011101100100: dataA <= 32'b01100010001001000000110110100001;
12'b011101100101: dataA <= 32'b00000110110101100010100101001111;
12'b011101100110: dataA <= 32'b01111100110000010101010010110000;
12'b011101100111: dataA <= 32'b00001001111110110001100111010010;
12'b011101101000: dataA <= 32'b10001000011010101101101100010010;
12'b011101101001: dataA <= 32'b00000110111110100011011000001010;
12'b011101101010: dataA <= 32'b11011110100000111010100110001011;
12'b011101101011: dataA <= 32'b00001011001111110010101100110110;
12'b011101101100: dataA <= 32'b00110110011010000101111001110011;
12'b011101101101: dataA <= 32'b00000110000111011110000110010111;
12'b011101101110: dataA <= 32'b10011100111001000111000101010101;
12'b011101101111: dataA <= 32'b00000111110111101110001101011100;
12'b011101110000: dataA <= 32'b11100110111010111101001110110001;
12'b011101110001: dataA <= 32'b00001011001000100111101010001100;
12'b011101110010: dataA <= 32'b00001001001111010100111111001110;
12'b011101110011: dataA <= 32'b00001000111110101100111000001011;
12'b011101110100: dataA <= 32'b10010011010100110101010110010001;
12'b011101110101: dataA <= 32'b00001001100001011101011001000001;
12'b011101110110: dataA <= 32'b10110111011010111111011111001101;
12'b011101110111: dataA <= 32'b00001000110111100101111011000110;
12'b011101111000: dataA <= 32'b01100000010110101101101110011000;
12'b011101111001: dataA <= 32'b00001001010101110000101101100000;
12'b011101111010: dataA <= 32'b00011000101110000011110111110110;
12'b011101111011: dataA <= 32'b00000111111110101110010001010100;
12'b011101111100: dataA <= 32'b10110100010100010101110010111011;
12'b011101111101: dataA <= 32'b00001000110100100011100110100101;
12'b011101111110: dataA <= 32'b01010110011010011010101000010111;
12'b011101111111: dataA <= 32'b00001101100110111100110100100001;
12'b011110000000: dataA <= 32'b11010010111001100110001010000011;
12'b011110000001: dataA <= 32'b00000100011101011110111001010001;
12'b011110000010: dataA <= 32'b11000110011100100110010011110100;
12'b011110000011: dataA <= 32'b00000011011000010011000100001100;
12'b011110000100: dataA <= 32'b11011000000101000000110110010101;
12'b011110000101: dataA <= 32'b00001010011010101101011000101011;
12'b011110000110: dataA <= 32'b00010011000101101011010110110010;
12'b011110000111: dataA <= 32'b00000101000110011100110000101011;
12'b011110001000: dataA <= 32'b10110001011101110111101011101001;
12'b011110001001: dataA <= 32'b00000010000110010000110011000100;
12'b011110001010: dataA <= 32'b11101110100101101111101000110000;
12'b011110001011: dataA <= 32'b00000010011001010110100010100100;
12'b011110001100: dataA <= 32'b01100010100011000100101101101000;
12'b011110001101: dataA <= 32'b00000011101110010100101001111011;
12'b011110001110: dataA <= 32'b00010011001100101110110101110101;
12'b011110001111: dataA <= 32'b00000101110111100010110000100101;
12'b011110010000: dataA <= 32'b10010111001101011001010100011001;
12'b011110010001: dataA <= 32'b00001010111010111010111101100001;
12'b011110010010: dataA <= 32'b11110101100110001111101010010111;
12'b011110010011: dataA <= 32'b00000101011000100010011010101011;
12'b011110010100: dataA <= 32'b00010110111110001010101010100100;
12'b011110010101: dataA <= 32'b00001010001100110000100000110100;
12'b011110010110: dataA <= 32'b11010010111011010011011100111011;
12'b011110010111: dataA <= 32'b00000011110011010110011000110100;
12'b011110011000: dataA <= 32'b10001110100001010101110110010011;
12'b011110011001: dataA <= 32'b00001001111000101110110000001011;
12'b011110011010: dataA <= 32'b10110101001111001010011110101001;
12'b011110011011: dataA <= 32'b00000001110100011000101111011011;
12'b011110011100: dataA <= 32'b00100001100110110111011101010000;
12'b011110011101: dataA <= 32'b00000110010001011100110010101001;
12'b011110011110: dataA <= 32'b00010110101110001110011100000111;
12'b011110011111: dataA <= 32'b00001001110110110001110000111110;
12'b011110100000: dataA <= 32'b00101101001010011011101011001001;
12'b011110100001: dataA <= 32'b00001101100110111000100010011110;
12'b011110100010: dataA <= 32'b10011011010010100110111101011010;
12'b011110100011: dataA <= 32'b00000101000001011110111101110000;
12'b011110100100: dataA <= 32'b10100110011010101100111100101111;
12'b011110100101: dataA <= 32'b00001101001000111001010001010111;
12'b011110100110: dataA <= 32'b10110110101110110010101110001001;
12'b011110100111: dataA <= 32'b00000011010010011010100111011001;
12'b011110101000: dataA <= 32'b00101011101101011011010111100010;
12'b011110101001: dataA <= 32'b00000111100110011111001010010101;
12'b011110101010: dataA <= 32'b00110100010100010101110110000001;
12'b011110101011: dataA <= 32'b00000101110101011011000110111011;
12'b011110101100: dataA <= 32'b01101000001110000110011010101000;
12'b011110101101: dataA <= 32'b00001000110100101000101001111101;
12'b011110101110: dataA <= 32'b11011010111001010000100110000101;
12'b011110101111: dataA <= 32'b00000000101111001010101100101110;
12'b011110110000: dataA <= 32'b00110101101010111100111101101101;
12'b011110110001: dataA <= 32'b00001110000111101101110111010101;
12'b011110110010: dataA <= 32'b00111100111010110011101011011010;
12'b011110110011: dataA <= 32'b00000010110111011010010111000100;
12'b011110110100: dataA <= 32'b11011010111100101001010011001001;
12'b011110110101: dataA <= 32'b00000110111001011111010001011100;
12'b011110110110: dataA <= 32'b01010100101001001001110010110110;
12'b011110110111: dataA <= 32'b00001011011011110001011001101000;
12'b011110111000: dataA <= 32'b00000000000010011001011001001010;
12'b011110111001: dataA <= 32'b00000000000000000000000000000000;
12'b011110111010: dataA <= 32'b10011110001000101001010101100001;
12'b011110111011: dataA <= 32'b00000111010101011110100001100111;
12'b011110111100: dataA <= 32'b11111010100100100101110010110011;
12'b011110111101: dataA <= 32'b00001011011101110101100011000001;
12'b011110111110: dataA <= 32'b01000100100110110101011100010000;
12'b011110111111: dataA <= 32'b00001000011110100101011000001011;
12'b011111000000: dataA <= 32'b01011010100000110011000101101100;
12'b011111000001: dataA <= 32'b00001011001110110000100101001111;
12'b011111000010: dataA <= 32'b11110010010010010101111001110010;
12'b011111000011: dataA <= 32'b00000101001000011000000110100110;
12'b011111000100: dataA <= 32'b11011100111001010111100101110110;
12'b011111000101: dataA <= 32'b00001000110111101010000101011100;
12'b011111000110: dataA <= 32'b11100110111010111100101110101111;
12'b011111000111: dataA <= 32'b00001010000111101011100110001100;
12'b011111001000: dataA <= 32'b11001011010111010100011110101011;
12'b011111001001: dataA <= 32'b00001010011110101100110100001011;
12'b011111001010: dataA <= 32'b00010101011001000101110110010010;
12'b011111001011: dataA <= 32'b00001000000001100001011100110010;
12'b011111001100: dataA <= 32'b01111001010011001110111110101010;
12'b011111001101: dataA <= 32'b00001001110111101001111011010110;
12'b011111001110: dataA <= 32'b10011010010110110101011110110110;
12'b011111001111: dataA <= 32'b00001001110101101110100101001000;
12'b011111010000: dataA <= 32'b01010110110010000011111000010110;
12'b011111010001: dataA <= 32'b00001001011110101010001101010100;
12'b011111010010: dataA <= 32'b01110000001100100110010100011100;
12'b011111010011: dataA <= 32'b00001001010100100111100110101101;
12'b011111010100: dataA <= 32'b00010010011110010010101001010111;
12'b011111010101: dataA <= 32'b00001101000100111010101000011010;
12'b011111010110: dataA <= 32'b01010001000001110110001001000011;
12'b011111010111: dataA <= 32'b00000101111110011110111001000010;
12'b011111011000: dataA <= 32'b10000100100100110110110100010110;
12'b011111011001: dataA <= 32'b00000011111010010011001000010101;
12'b011111011010: dataA <= 32'b10010010001000101001010110110101;
12'b011111011011: dataA <= 32'b00001011011001101111010000101100;
12'b011111011100: dataA <= 32'b10010011001001101011010110110010;
12'b011111011101: dataA <= 32'b00000100000111011010110000101011;
12'b011111011110: dataA <= 32'b00110011010110001111101010101000;
12'b011111011111: dataA <= 32'b00000001001001010000111011000100;
12'b011111100000: dataA <= 32'b10101010100010000111101000110000;
12'b011111100001: dataA <= 32'b00000011011011010010100110100100;
12'b011111100010: dataA <= 32'b01011110011111000100001101000101;
12'b011111100011: dataA <= 32'b00000011010000010010101101111011;
12'b011111100100: dataA <= 32'b10010101010001000111000110010110;
12'b011111100101: dataA <= 32'b00000110110111100000110000101101;
12'b011111100110: dataA <= 32'b11011001010001001001100100111010;
12'b011111100111: dataA <= 32'b00001011111001111010110101010001;
12'b011111101000: dataA <= 32'b10111001011110100111101011010110;
12'b011111101001: dataA <= 32'b00000110011001011110010110101011;
12'b011111101010: dataA <= 32'b10010111000010000010101001100011;
12'b011111101011: dataA <= 32'b00001001101011101100011000110100;
12'b011111101100: dataA <= 32'b01010001000011001010111101111001;
12'b011111101101: dataA <= 32'b00000100010101010010011100111101;
12'b011111101110: dataA <= 32'b01001100101001100110000110110011;
12'b011111101111: dataA <= 32'b00001010110111101100101100001100;
12'b011111110000: dataA <= 32'b00110101000110111001111110000111;
12'b011111110001: dataA <= 32'b00000010010110010110110011010011;
12'b011111110010: dataA <= 32'b11100101100111000110111101001110;
12'b011111110011: dataA <= 32'b00000110010001011100110010011000;
12'b011111110100: dataA <= 32'b10010100110010011110011011100101;
12'b011111110101: dataA <= 32'b00001010010101110101101001000110;
12'b011111110110: dataA <= 32'b11101101000110011011101010001000;
12'b011111110111: dataA <= 32'b00001100100100110100010110101101;
12'b011111111000: dataA <= 32'b10011101010010110110101110011000;
12'b011111111001: dataA <= 32'b00000100000011011110111101100000;
12'b011111111010: dataA <= 32'b10100010011010101100101100101101;
12'b011111111011: dataA <= 32'b00001100000110111001001001101111;
12'b011111111100: dataA <= 32'b00110100100110101010011101000111;
12'b011111111101: dataA <= 32'b00000011110100011000100111001001;
12'b011111111110: dataA <= 32'b11110001100101011011100110100010;
12'b011111111111: dataA <= 32'b00000110100110011111001010011100;
12'b100000000000: dataA <= 32'b11110000001100100110010100100010;
12'b100000000001: dataA <= 32'b00000110010110011011000110110010;
12'b100000000010: dataA <= 32'b01100100001110010110011001100111;
12'b100000000011: dataA <= 32'b00001001010100100110100110000101;
12'b100000000100: dataA <= 32'b00011010111000111000110101000110;
12'b100000000101: dataA <= 32'b00000000110010001010110101000111;
12'b100000000110: dataA <= 32'b10111001100010111100011101001011;
12'b100000000111: dataA <= 32'b00001101000101110001110011010100;
12'b100000001000: dataA <= 32'b10111010101110110011011100011000;
12'b100000001001: dataA <= 32'b00000011111001010110011011000011;
12'b100000001010: dataA <= 32'b00011010111100011001110010101011;
12'b100000001011: dataA <= 32'b00000111111001100001010001100101;
12'b100000001100: dataA <= 32'b10010010101100111010010011111000;
12'b100000001101: dataA <= 32'b00001100111001110011010001010000;
12'b100000001110: dataA <= 32'b00000000000010001001011000101010;
12'b100000001111: dataA <= 32'b00000000000000000000000000000000;
12'b100000010000: dataA <= 32'b11000101000000101110100000110100;
12'b100000010001: dataA <= 32'b00001010110001010001000011110100;
12'b100000010010: dataA <= 32'b11010010001010111110111001111010;
12'b100000010011: dataA <= 32'b00001110101001110000010100111001;
12'b100000010100: dataA <= 32'b10010011110110101010011000000111;
12'b100000010101: dataA <= 32'b00001111001111101100110101101111;
12'b100000010110: dataA <= 32'b10010001001001100110010110010100;
12'b100000010111: dataA <= 32'b00000111001001010010011111101101;
12'b100000011000: dataA <= 32'b11001000011010111011011001001100;
12'b100000011001: dataA <= 32'b00000100010101000011001111011010;
12'b100000011010: dataA <= 32'b00011101000111110101011011010100;
12'b100000011011: dataA <= 32'b00001011101110000010101010011101;
12'b100000011100: dataA <= 32'b10011100110010010010000111100010;
12'b100000011101: dataA <= 32'b00000011101011110010101010011011;
12'b100000011110: dataA <= 32'b10101011101010001001010101100010;
12'b100000011111: dataA <= 32'b00001111001011011010100101111111;
12'b100000100000: dataA <= 32'b01101101010110111101111001010011;
12'b100000100001: dataA <= 32'b00000000101111101110111101000110;
12'b100000100010: dataA <= 32'b01101000001111011001100101000010;
12'b100000100011: dataA <= 32'b00001011101100111100101111001001;
12'b100000100100: dataA <= 32'b10001011001010101010011011000010;
12'b100000100101: dataA <= 32'b00001010101100010010100000010101;
12'b100000100110: dataA <= 32'b01011001010001111011111011001111;
12'b100000100111: dataA <= 32'b00001111001101000110101010001101;
12'b100000101000: dataA <= 32'b10000110011111001110111110010111;
12'b100000101001: dataA <= 32'b00001010001101110010110010101010;
12'b100000101010: dataA <= 32'b00001111011001010011011011101101;
12'b100000101011: dataA <= 32'b00000010000101010100001001000111;
12'b100000101100: dataA <= 32'b11100001011111000100010001101101;
12'b100000101101: dataA <= 32'b00001111010100011101000001001101;
12'b100000101110: dataA <= 32'b01010011110111011110011011010111;
12'b100000101111: dataA <= 32'b00001101011000100101011010110111;
12'b100000110000: dataA <= 32'b10000101011000101110101010110010;
12'b100000110001: dataA <= 32'b00001100101001101000100010010110;
12'b100000110010: dataA <= 32'b10100101011001101100101001010010;
12'b100000110011: dataA <= 32'b00000011110111011001001001110110;
12'b100000110100: dataA <= 32'b11101010011011110011100100001010;
12'b100000110101: dataA <= 32'b00000100111101011101011110000001;
12'b100000110110: dataA <= 32'b11010000101011110011111000001110;
12'b100000110111: dataA <= 32'b00001101111001010011011010010010;
12'b100000111000: dataA <= 32'b00001111000010000001110010100101;
12'b100000111001: dataA <= 32'b00001000011001010111011001101100;
12'b100000111010: dataA <= 32'b10101001010111100101111011010011;
12'b100000111011: dataA <= 32'b00001011110010011000111110110110;
12'b100000111100: dataA <= 32'b01101001001100110101101101010110;
12'b100000111101: dataA <= 32'b00001100101000011010001000111101;
12'b100000111110: dataA <= 32'b10101110001111110010111011001001;
12'b100000111111: dataA <= 32'b00001100110011001011000001110010;
12'b100001000000: dataA <= 32'b01100001010001010011110001101100;
12'b100001000001: dataA <= 32'b00000101101100001100100110010110;
12'b100001000010: dataA <= 32'b00100001011101011001101100100100;
12'b100001000011: dataA <= 32'b00001010110111001111011010101110;
12'b100001000100: dataA <= 32'b10010101100111000100111001110010;
12'b100001000101: dataA <= 32'b00001011101010010110100110001111;
12'b100001000110: dataA <= 32'b01100010010100111010000011100011;
12'b100001000111: dataA <= 32'b00001011011011011001010001100001;
12'b100001001000: dataA <= 32'b00110010110111011001110111000101;
12'b100001001001: dataA <= 32'b00001000110011011001000100011011;
12'b100001001010: dataA <= 32'b11011001010111001011000010101000;
12'b100001001011: dataA <= 32'b00001010101011110100010111010101;
12'b100001001100: dataA <= 32'b10100010100101110011000100001011;
12'b100001001101: dataA <= 32'b00000010000110001010010110111010;
12'b100001001110: dataA <= 32'b11101001000111010010011100000011;
12'b100001001111: dataA <= 32'b00000001110111011111000000010100;
12'b100001010000: dataA <= 32'b10001100111010010010100110100110;
12'b100001010001: dataA <= 32'b00000011000111100100001111110100;
12'b100001010010: dataA <= 32'b10010010010101001010100011100101;
12'b100001010011: dataA <= 32'b00001010011000010011001100100001;
12'b100001010100: dataA <= 32'b00110010011101110101000001010010;
12'b100001010101: dataA <= 32'b00000011010010100101000010011011;
12'b100001010110: dataA <= 32'b01000110011111001110110001010110;
12'b100001010111: dataA <= 32'b00001011010011100011001001011010;
12'b100001011000: dataA <= 32'b11000110110111001011010011101100;
12'b100001011001: dataA <= 32'b00001010001101010010110010101011;
12'b100001011010: dataA <= 32'b11011101001000011110000011010101;
12'b100001011011: dataA <= 32'b00001001011110011011101011100101;
12'b100001011100: dataA <= 32'b01110000001110001010000101100101;
12'b100001011101: dataA <= 32'b00000010100101111000011110010001;
12'b100001011110: dataA <= 32'b11010110001001101010011100000111;
12'b100001011111: dataA <= 32'b00001100111000001101010001110001;
12'b100001100000: dataA <= 32'b11011111001000111111000101111010;
12'b100001100001: dataA <= 32'b00001100110000101000111110100100;
12'b100001100010: dataA <= 32'b01010111011001001110001100011000;
12'b100001100011: dataA <= 32'b00001100100110101000011000010101;
12'b100001100100: dataA <= 32'b00000000000000101011100101001110;
12'b100001100101: dataA <= 32'b00000000000000000000000000000000;
12'b100001100110: dataA <= 32'b10000100111000011101110000110010;
12'b100001100111: dataA <= 32'b00001010110010010010111011101101;
12'b100001101000: dataA <= 32'b01011000000110101111011000011010;
12'b100001101001: dataA <= 32'b00001111001100110010011101001001;
12'b100001101010: dataA <= 32'b10001101101110110010101001000111;
12'b100001101011: dataA <= 32'b00001111010010101100111001010111;
12'b100001101100: dataA <= 32'b01010001000001010110000101110011;
12'b100001101101: dataA <= 32'b00000111101001010110011011011110;
12'b100001101110: dataA <= 32'b01001100010010111011111001101100;
12'b100001101111: dataA <= 32'b00000011110011000011000011100011;
12'b100001110000: dataA <= 32'b00011101000111100101111010110101;
12'b100001110001: dataA <= 32'b00001011110000000110100010010101;
12'b100001110010: dataA <= 32'b10011100110010100010001000100010;
12'b100001110011: dataA <= 32'b00000100001001110100110010011011;
12'b100001110100: dataA <= 32'b10100111101110011001010111000001;
12'b100001110101: dataA <= 32'b00001111001110011100100101100111;
12'b100001110110: dataA <= 32'b11101011011010101110011000110011;
12'b100001110111: dataA <= 32'b00000000101100101101000100110101;
12'b100001111000: dataA <= 32'b11101100010011101010000110100001;
12'b100001111001: dataA <= 32'b00001011101110111100110111010001;
12'b100001111010: dataA <= 32'b11001010111110110010101100000011;
12'b100001111011: dataA <= 32'b00001010101101010110011100001100;
12'b100001111100: dataA <= 32'b01010111001101111011111011010000;
12'b100001111101: dataA <= 32'b00001111010000001000100010000101;
12'b100001111110: dataA <= 32'b11001010010110111111011101111010;
12'b100001111111: dataA <= 32'b00001010001110110010111010110010;
12'b100010000000: dataA <= 32'b11001101010001010011001011101111;
12'b100010000001: dataA <= 32'b00000011000100011010000100101110;
12'b100010000010: dataA <= 32'b01011101011011000100110001101011;
12'b100010000011: dataA <= 32'b00001110110111011101000000111101;
12'b100010000100: dataA <= 32'b10001111110011001110111010011000;
12'b100010000101: dataA <= 32'b00001100011001100011011010011111;
12'b100010000110: dataA <= 32'b10000011001100011101111010110011;
12'b100010000111: dataA <= 32'b00001101001011101100100101111110;
12'b100010001000: dataA <= 32'b10100011011001101100101001010010;
12'b100010001001: dataA <= 32'b00000011010101011001000101100110;
12'b100010001010: dataA <= 32'b11101110011111110100010100101000;
12'b100010001011: dataA <= 32'b00000011011011011001011110010001;
12'b100010001100: dataA <= 32'b11010010100011110100101000001110;
12'b100010001101: dataA <= 32'b00001100111011010001010010011010;
12'b100010001110: dataA <= 32'b00010000111010010001110100000100;
12'b100010001111: dataA <= 32'b00000111011000010101010101101100;
12'b100010010000: dataA <= 32'b11100111011011011110101010110100;
12'b100010010001: dataA <= 32'b00001011110100011000111010100110;
12'b100010010010: dataA <= 32'b11100111010000101101001100110111;
12'b100010010011: dataA <= 32'b00001101001010011110001000110100;
12'b100010010100: dataA <= 32'b10110010010111110011101011101011;
12'b100010010101: dataA <= 32'b00001100010101001100111001111010;
12'b100010010110: dataA <= 32'b01011111010001010011100010001010;
12'b100010010111: dataA <= 32'b00000110001011010000011110000110;
12'b100010011000: dataA <= 32'b01011101011001101001011101100110;
12'b100010011001: dataA <= 32'b00001001111000001101010010011110;
12'b100010011010: dataA <= 32'b10010001100010111101011001110011;
12'b100010011011: dataA <= 32'b00001100001100011000100001110111;
12'b100010011100: dataA <= 32'b00100110010101001001100100100010;
12'b100010011101: dataA <= 32'b00001010011100010111001101110001;
12'b100010011110: dataA <= 32'b10110010111111101010011000000101;
12'b100010011111: dataA <= 32'b00001000110011011001000100100010;
12'b100010100000: dataA <= 32'b00010111010011001011100011100111;
12'b100010100001: dataA <= 32'b00001011001100111000011111000110;
12'b100010100010: dataA <= 32'b00100100100101110011000100101001;
12'b100010100011: dataA <= 32'b00000011000100010000001111000011;
12'b100010100100: dataA <= 32'b01101001001011011010111101000101;
12'b100010100101: dataA <= 32'b00000000110101011111000000010100;
12'b100010100110: dataA <= 32'b01001100110010011010100111100110;
12'b100010100111: dataA <= 32'b00000100000101101000001111110101;
12'b100010101000: dataA <= 32'b00010110010001010010010100100011;
12'b100010101001: dataA <= 32'b00001001011001010011001000110001;
12'b100010101010: dataA <= 32'b01110110101001101101000001010000;
12'b100010101011: dataA <= 32'b00000011010000100101000010100011;
12'b100010101100: dataA <= 32'b00001010010110111111010000110011;
12'b100010101101: dataA <= 32'b00001010110100100011001001100010;
12'b100010101110: dataA <= 32'b00000110101111001011110100001010;
12'b100010101111: dataA <= 32'b00001010001110010100101110101100;
12'b100010110000: dataA <= 32'b10011101001000010101010010110011;
12'b100010110001: dataA <= 32'b00000111111110010111101011011110;
12'b100010110010: dataA <= 32'b01110100010110011010000110100100;
12'b100010110011: dataA <= 32'b00000011100011111010100110100001;
12'b100010110100: dataA <= 32'b11011100000101110010011101001001;
12'b100010110101: dataA <= 32'b00001011111010001011001010000001;
12'b100010110110: dataA <= 32'b00011111001000101110100100111001;
12'b100010110111: dataA <= 32'b00001100110010101001000010011101;
12'b100010111000: dataA <= 32'b10010101010100111101101011011010;
12'b100010111001: dataA <= 32'b00001101101001101100011100001100;
12'b100010111010: dataA <= 32'b00000000000000101011000101001101;
12'b100010111011: dataA <= 32'b00000000000000000000000000000000;
12'b100010111100: dataA <= 32'b00000110101100001101010000101111;
12'b100010111101: dataA <= 32'b00001010010011010010110111100110;
12'b100010111110: dataA <= 32'b00011110000110010111010111011010;
12'b100010111111: dataA <= 32'b00001111001111110110100101011001;
12'b100011000000: dataA <= 32'b00001001100110111011001010001000;
12'b100011000001: dataA <= 32'b00001111010101101101000001000111;
12'b100011000010: dataA <= 32'b11010000111101000101110101010010;
12'b100011000011: dataA <= 32'b00001000101001011010010111001110;
12'b100011000100: dataA <= 32'b11010000001010111100001001101101;
12'b100011000101: dataA <= 32'b00000011010001000010110111100011;
12'b100011000110: dataA <= 32'b01011101000111010110101010010110;
12'b100011000111: dataA <= 32'b00001011110001001010010110001101;
12'b100011001000: dataA <= 32'b11011110110010101010011010000011;
12'b100011001001: dataA <= 32'b00000100101000110100111010011011;
12'b100011001010: dataA <= 32'b01100011110010101001101000000001;
12'b100011001011: dataA <= 32'b00001111010001100000100101001111;
12'b100011001100: dataA <= 32'b01100111011110011110011000110100;
12'b100011001101: dataA <= 32'b00000001001001101101001000101101;
12'b100011001110: dataA <= 32'b10110000010111110010110111100001;
12'b100011001111: dataA <= 32'b00001100001111111101000011100010;
12'b100011010000: dataA <= 32'b00001010110110111011001101000101;
12'b100011010001: dataA <= 32'b00001011001110011010011000001100;
12'b100011010010: dataA <= 32'b01010101001001111011111010110001;
12'b100011010011: dataA <= 32'b00001111010011001100011001111101;
12'b100011010100: dataA <= 32'b01001110001110100111101100011100;
12'b100011010101: dataA <= 32'b00001010001111110011000010111011;
12'b100011010110: dataA <= 32'b00001011001001011010111011110000;
12'b100011010111: dataA <= 32'b00000100100010011110000100011110;
12'b100011011000: dataA <= 32'b00011011011010111101010010101000;
12'b100011011001: dataA <= 32'b00001101111001011101000000110101;
12'b100011011010: dataA <= 32'b10001011101010111111011001011001;
12'b100011011011: dataA <= 32'b00001011011011011111011010000111;
12'b100011011100: dataA <= 32'b10000011000000001101011010010100;
12'b100011011101: dataA <= 32'b00001101101110101110101001101110;
12'b100011011110: dataA <= 32'b01011111011001100100011000110011;
12'b100011011111: dataA <= 32'b00000010110011010111000101010110;
12'b100011100000: dataA <= 32'b00110010100111110101000101100111;
12'b100011100001: dataA <= 32'b00000010011001010111011010100010;
12'b100011100010: dataA <= 32'b00010110011111110101011000001110;
12'b100011100011: dataA <= 32'b00001011111101001111001110100011;
12'b100011100100: dataA <= 32'b11010000110110100010000101000010;
12'b100011100101: dataA <= 32'b00000110011000010011010001101011;
12'b100011100110: dataA <= 32'b00100101011011000111001010010101;
12'b100011100111: dataA <= 32'b00001011010101011000111010010111;
12'b100011101000: dataA <= 32'b01100101010100100100011011111001;
12'b100011101001: dataA <= 32'b00001101101101100100001000110100;
12'b100011101010: dataA <= 32'b10110110011111110100011100001100;
12'b100011101011: dataA <= 32'b00001011110111001100110010000010;
12'b100011101100: dataA <= 32'b01011101001101010011010010101000;
12'b100011101101: dataA <= 32'b00000110101010010100010101110110;
12'b100011101110: dataA <= 32'b01011011011001111001011110101001;
12'b100011101111: dataA <= 32'b00001000111001001011001010001110;
12'b100011110000: dataA <= 32'b10001101011010110101101001010011;
12'b100011110001: dataA <= 32'b00001100101110011100100001011111;
12'b100011110010: dataA <= 32'b00101010011001011001010110000001;
12'b100011110011: dataA <= 32'b00001000111101010101001010000001;
12'b100011110100: dataA <= 32'b00110011000111110011001001000110;
12'b100011110101: dataA <= 32'b00001000010011011001000000101010;
12'b100011110110: dataA <= 32'b10010101001111001100000100100101;
12'b100011110111: dataA <= 32'b00001011001101111010101010110110;
12'b100011111000: dataA <= 32'b10101000101001111011000101001000;
12'b100011111001: dataA <= 32'b00000100000011010100000111001011;
12'b100011111010: dataA <= 32'b10100111001111100011011110000111;
12'b100011111011: dataA <= 32'b00000000110010011111000000010011;
12'b100011111100: dataA <= 32'b11001110101010100010111000100110;
12'b100011111101: dataA <= 32'b00000101000100101110010111100101;
12'b100011111110: dataA <= 32'b11011010001101100010000101100010;
12'b100011111111: dataA <= 32'b00001000011001010001000001000000;
12'b100100000000: dataA <= 32'b01111000110001100100110001001101;
12'b100100000001: dataA <= 32'b00000011001110100101000110100011;
12'b100100000010: dataA <= 32'b00001110001110100111100000110000;
12'b100100000011: dataA <= 32'b00001010010101100001001001110010;
12'b100100000100: dataA <= 32'b01001010100011001100010100101001;
12'b100100000101: dataA <= 32'b00001010001111010110101010100100;
12'b100100000110: dataA <= 32'b00011011001000001100110010110001;
12'b100100000111: dataA <= 32'b00000110011110010011100111000111;
12'b100100001000: dataA <= 32'b10111000011110100010010111100100;
12'b100100001001: dataA <= 32'b00000101000010111100110010110001;
12'b100100001010: dataA <= 32'b00100000000110000010011101101011;
12'b100100001011: dataA <= 32'b00001010111011001011000010010010;
12'b100100001100: dataA <= 32'b01011101001000011110000100011000;
12'b100100001101: dataA <= 32'b00001100010100100111000110010101;
12'b100100001110: dataA <= 32'b11010011010000110101011010011011;
12'b100100001111: dataA <= 32'b00001110001011110000100100001011;
12'b100100010000: dataA <= 32'b00000000000000110010100101101100;
12'b100100010001: dataA <= 32'b00000000000000000000000000000000;
12'b100100010010: dataA <= 32'b10001000100100001100100000101100;
12'b100100010011: dataA <= 32'b00001010010100010010110011010110;
12'b100100010100: dataA <= 32'b00100100000101111111100110011010;
12'b100100010101: dataA <= 32'b00001111010010111000101101110001;
12'b100100010110: dataA <= 32'b10000101011111000011011010101001;
12'b100100010111: dataA <= 32'b00001110010111101101000100101110;
12'b100100011000: dataA <= 32'b01010000110100111101010101010001;
12'b100100011001: dataA <= 32'b00001001001010011110010110111111;
12'b100100011010: dataA <= 32'b10010110000110111100101010001110;
12'b100100011011: dataA <= 32'b00000011010000000010101011100100;
12'b100100011100: dataA <= 32'b01011011000011000111001001010111;
12'b100100011101: dataA <= 32'b00001011010010001110001110000101;
12'b100100011110: dataA <= 32'b00100000110010110010111011000100;
12'b100100011111: dataA <= 32'b00000101100111110101000110011100;
12'b100100100000: dataA <= 32'b00011111110010110001111001100010;
12'b100100100001: dataA <= 32'b00001111010100100010100100111111;
12'b100100100010: dataA <= 32'b11100101100010001110101000010100;
12'b100100100011: dataA <= 32'b00000001100111101101001100100100;
12'b100100100100: dataA <= 32'b00110100011111110011101001000001;
12'b100100100101: dataA <= 32'b00001011110001111101001111101011;
12'b100100100110: dataA <= 32'b01001100101111000011011110001000;
12'b100100100111: dataA <= 32'b00001011010000011110011000001011;
12'b100100101000: dataA <= 32'b01010101000101111011111010110011;
12'b100100101001: dataA <= 32'b00001110110110010000010001110101;
12'b100100101010: dataA <= 32'b10010100001010001111101011011101;
12'b100100101011: dataA <= 32'b00001010010000110011001010111011;
12'b100100101100: dataA <= 32'b10001011000001100010101011110010;
12'b100100101101: dataA <= 32'b00000110000001100100000100010101;
12'b100100101110: dataA <= 32'b10011001011010110101100011000110;
12'b100100101111: dataA <= 32'b00001100111011011101000000110100;
12'b100100110000: dataA <= 32'b10000111011110100111101000011001;
12'b100100110001: dataA <= 32'b00001010011100011101011001101111;
12'b100100110010: dataA <= 32'b01000010110100001100101001110101;
12'b100100110011: dataA <= 32'b00001101110000110000110001011110;
12'b100100110100: dataA <= 32'b00011101011001100100011000110011;
12'b100100110101: dataA <= 32'b00000010010001010111000001001110;
12'b100100110110: dataA <= 32'b01110100101111101101110110000111;
12'b100100110111: dataA <= 32'b00000001010111010101010110101010;
12'b100100111000: dataA <= 32'b01011000011111100101111000101110;
12'b100100111001: dataA <= 32'b00001010011110001101000110100011;
12'b100100111010: dataA <= 32'b11010010101110101010010110100010;
12'b100100111011: dataA <= 32'b00000101110111010001001001101011;
12'b100100111100: dataA <= 32'b00100001011110110111011001110110;
12'b100100111101: dataA <= 32'b00001010010110011000110101111111;
12'b100100111110: dataA <= 32'b11100011010100100011111010111010;
12'b100100111111: dataA <= 32'b00001110001111101010001100110011;
12'b100101000000: dataA <= 32'b10111000100111110101001100101110;
12'b100101000001: dataA <= 32'b00001010111000001110101010001010;
12'b100101000010: dataA <= 32'b00011101001101011011000011100110;
12'b100101000011: dataA <= 32'b00000111001010011000010101100110;
12'b100101000100: dataA <= 32'b01011001011010001001011111001011;
12'b100101000101: dataA <= 32'b00001000011001001011000001111110;
12'b100101000110: dataA <= 32'b01001011010010101110001000110100;
12'b100101000111: dataA <= 32'b00001100101111011110100001000111;
12'b100101001000: dataA <= 32'b01101100011101101001000111100001;
12'b100101001001: dataA <= 32'b00000111111101010101000110010001;
12'b100101001010: dataA <= 32'b10110001001111110011111010000111;
12'b100101001011: dataA <= 32'b00000111110011011000111100111001;
12'b100101001100: dataA <= 32'b11010011001011001100100101100100;
12'b100101001101: dataA <= 32'b00001011101111111100110110100110;
12'b100101001110: dataA <= 32'b11101010101110000011000110000111;
12'b100101001111: dataA <= 32'b00000101100001011010000111001011;
12'b100101010000: dataA <= 32'b11100111001111100100001110101010;
12'b100101010001: dataA <= 32'b00000000101111011111000000010010;
12'b100101010010: dataA <= 32'b10010000100010101011001001100111;
12'b100101010011: dataA <= 32'b00000110100011110010011011010110;
12'b100101010100: dataA <= 32'b01100000001101101001110111000001;
12'b100101010101: dataA <= 32'b00000111011001010000111101011000;
12'b100101010110: dataA <= 32'b10111000111001100100110001101010;
12'b100101010111: dataA <= 32'b00000011101100100101000110100011;
12'b100101011000: dataA <= 32'b00010100001010001111100000101101;
12'b100101011001: dataA <= 32'b00001001110110100001001001111010;
12'b100101011010: dataA <= 32'b10001100011011000100110101000111;
12'b100101011011: dataA <= 32'b00001010010000011000100110100100;
12'b100101011100: dataA <= 32'b01011011000100001100000010101110;
12'b100101011101: dataA <= 32'b00000100111101010001011110110111;
12'b100101011110: dataA <= 32'b00111010101010101010101000100100;
12'b100101011111: dataA <= 32'b00000110100001111100111110111010;
12'b100101100000: dataA <= 32'b00100110001010001010011101101110;
12'b100101100001: dataA <= 32'b00001001011100001010111010011010;
12'b100101100010: dataA <= 32'b01011101001000010101010011010110;
12'b100101100011: dataA <= 32'b00001011110110100111000110001101;
12'b100101100100: dataA <= 32'b01010001001000101100111000111011;
12'b100101100101: dataA <= 32'b00001110101101110010101000001011;
12'b100101100110: dataA <= 32'b00000000000000111010010101101011;
12'b100101100111: dataA <= 32'b00000000000000000000000000000000;
12'b100101101000: dataA <= 32'b00001100011100001011110001001001;
12'b100101101001: dataA <= 32'b00001001110101010100101110111111;
12'b100101101010: dataA <= 32'b11101000000101101111010101011001;
12'b100101101011: dataA <= 32'b00001111010101111000111010000000;
12'b100101101100: dataA <= 32'b00000011010011000011111011001010;
12'b100101101101: dataA <= 32'b00001101011010101101001000011110;
12'b100101101110: dataA <= 32'b10010010110000110101000101010000;
12'b100101101111: dataA <= 32'b00001001101010100010010110100111;
12'b100101110000: dataA <= 32'b00011100000110110100111010001111;
12'b100101110001: dataA <= 32'b00000011001110000110100011011101;
12'b100101110010: dataA <= 32'b01011011000010110111011000110111;
12'b100101110011: dataA <= 32'b00001010110100010010001001111101;
12'b100101110100: dataA <= 32'b01100010110010111011001100000110;
12'b100101110101: dataA <= 32'b00000110100110110101001110011100;
12'b100101110110: dataA <= 32'b10011001101111000010011011000011;
12'b100101110111: dataA <= 32'b00001110110111100100100100101110;
12'b100101111000: dataA <= 32'b00100001100001111110100111110100;
12'b100101111001: dataA <= 32'b00000010100101101011010000011100;
12'b100101111010: dataA <= 32'b11110110101011110100011010100010;
12'b100101111011: dataA <= 32'b00001011110010111011011011101011;
12'b100101111100: dataA <= 32'b11001110101011000011111111001010;
12'b100101111101: dataA <= 32'b00001011010001100000011000001010;
12'b100101111110: dataA <= 32'b00010101000001111011111010010100;
12'b100101111111: dataA <= 32'b00001110011000010100001101101101;
12'b100110000000: dataA <= 32'b00011010000101110111101001111110;
12'b100110000001: dataA <= 32'b00001010010001110001010010111100;
12'b100110000010: dataA <= 32'b11001010111001101010101011010011;
12'b100110000011: dataA <= 32'b00000111100001101010001000001100;
12'b100110000100: dataA <= 32'b00010111010110100101110100000101;
12'b100110000101: dataA <= 32'b00001011111101011100111100110100;
12'b100110000110: dataA <= 32'b10000011010110001111100111111001;
12'b100110000111: dataA <= 32'b00001000111100011011011001010111;
12'b100110001000: dataA <= 32'b00000010101000001011111001010101;
12'b100110001001: dataA <= 32'b00001101110010110000111001010110;
12'b100110001010: dataA <= 32'b10011011011001100100001000010011;
12'b100110001011: dataA <= 32'b00000010001110010110111100111101;
12'b100110001100: dataA <= 32'b10110100110111011110010111000110;
12'b100110001101: dataA <= 32'b00000000110100010011010010110010;
12'b100110001110: dataA <= 32'b10011100011011010110101000101110;
12'b100110001111: dataA <= 32'b00001000111110001100111110101011;
12'b100110010000: dataA <= 32'b11010100101010110010100111100001;
12'b100110010001: dataA <= 32'b00000100110110010001000101101011;
12'b100110010010: dataA <= 32'b00011111011110011111101001010111;
12'b100110010011: dataA <= 32'b00001001110111011010110001101111;
12'b100110010100: dataA <= 32'b01100001010100100011011001111011;
12'b100110010101: dataA <= 32'b00001101110001101110010000110011;
12'b100110010110: dataA <= 32'b11111010110011101101111100110000;
12'b100110010111: dataA <= 32'b00001010011001010000100010010010;
12'b100110011000: dataA <= 32'b00011011001101100010110100100100;
12'b100110011001: dataA <= 32'b00000111101010011100010001010110;
12'b100110011010: dataA <= 32'b01010111010110011001101111001110;
12'b100110011011: dataA <= 32'b00000111011001001010111001101110;
12'b100110011100: dataA <= 32'b11001011001010011110001000010100;
12'b100110011101: dataA <= 32'b00001100110001100010100000110110;
12'b100110011110: dataA <= 32'b01110000100101111001001001000001;
12'b100110011111: dataA <= 32'b00000110011101010101000010100001;
12'b100110100000: dataA <= 32'b00110001010111110100101011001000;
12'b100110100001: dataA <= 32'b00000111010011011000111001001001;
12'b100110100010: dataA <= 32'b00010011000111000101000110100011;
12'b100110100011: dataA <= 32'b00001011110000111101000010010111;
12'b100110100100: dataA <= 32'b01101100110010001011000111000111;
12'b100110100101: dataA <= 32'b00000110100001100000000111001100;
12'b100110100110: dataA <= 32'b01100101010011100100101111001101;
12'b100110100111: dataA <= 32'b00000000101100011111000000011010;
12'b100110101000: dataA <= 32'b00010100011110101011011010100111;
12'b100110101001: dataA <= 32'b00000111100011110100100011000111;
12'b100110101010: dataA <= 32'b01100100001101111001111000100001;
12'b100110101011: dataA <= 32'b00000110011000010010110101101000;
12'b100110101100: dataA <= 32'b11111001000101011100100010001000;
12'b100110101101: dataA <= 32'b00000011101010100011001010100011;
12'b100110101110: dataA <= 32'b00011010000101110111100000101011;
12'b100110101111: dataA <= 32'b00001001010111011111001010001010;
12'b100110110000: dataA <= 32'b11010000010111000101010110000111;
12'b100110110001: dataA <= 32'b00001010010001011010100010011100;
12'b100110110010: dataA <= 32'b10011011000100001011010010101100;
12'b100110110011: dataA <= 32'b00000011111100001101011010011111;
12'b100110110100: dataA <= 32'b01111100110110110010111001100101;
12'b100110110101: dataA <= 32'b00001000000001111101001011001010;
12'b100110110110: dataA <= 32'b01101100001110010010011110010000;
12'b100110110111: dataA <= 32'b00001000011100001100110010100010;
12'b100110111000: dataA <= 32'b01011011000100001100100010110100;
12'b100110111001: dataA <= 32'b00001011010111100111001010000101;
12'b100110111010: dataA <= 32'b10010001000100101100010111111100;
12'b100110111011: dataA <= 32'b00001110110000110100110000010010;
12'b100110111100: dataA <= 32'b00000000000001001001110110001010;
12'b100110111101: dataA <= 32'b00000000000000000000000000000000;
12'b100110111110: dataA <= 32'b10010000010100001011000001100111;
12'b100110111111: dataA <= 32'b00001000110101010110101010101111;
12'b100111000000: dataA <= 32'b00101110001101010111010100111000;
12'b100111000001: dataA <= 32'b00001110010111111011000010010001;
12'b100111000010: dataA <= 32'b10000011000111000100011011101011;
12'b100111000011: dataA <= 32'b00001100011100101011001100010101;
12'b100111000100: dataA <= 32'b10010100101100101100100101001111;
12'b100111000101: dataA <= 32'b00001010001011100110011010001111;
12'b100111000110: dataA <= 32'b10100010000110101101001010001111;
12'b100111000111: dataA <= 32'b00000011101100001010010111010101;
12'b100111001000: dataA <= 32'b01011011000010011111100111111000;
12'b100111001001: dataA <= 32'b00001010110101011000000101110101;
12'b100111001010: dataA <= 32'b01100010110010111011011101001000;
12'b100111001011: dataA <= 32'b00000111100110110011010110011100;
12'b100111001100: dataA <= 32'b11010101101011001010101100000100;
12'b100111001101: dataA <= 32'b00001101111001100110101000011101;
12'b100111001110: dataA <= 32'b10011101100001101110100111010100;
12'b100111001111: dataA <= 32'b00000100000011101001010100011011;
12'b100111010000: dataA <= 32'b01111000110011110101001100000011;
12'b100111010001: dataA <= 32'b00001011010100111001100011101100;
12'b100111010010: dataA <= 32'b00010000100011000100011111001101;
12'b100111010011: dataA <= 32'b00001010110010100100011000011010;
12'b100111010100: dataA <= 32'b00010100111101111011111001110100;
12'b100111010101: dataA <= 32'b00001101011010011010001001100101;
12'b100111010110: dataA <= 32'b01100000000101011111101000011110;
12'b100111010111: dataA <= 32'b00001010010010101111011010111100;
12'b100111011000: dataA <= 32'b00001100110001110010011010110100;
12'b100111011001: dataA <= 32'b00001001000001110000001100001100;
12'b100111011010: dataA <= 32'b10010101010010011110000101000100;
12'b100111011011: dataA <= 32'b00001010011110011100111100110011;
12'b100111011100: dataA <= 32'b00000011001001110111100110111001;
12'b100111011101: dataA <= 32'b00000111111101011001010101000111;
12'b100111011110: dataA <= 32'b11000110100000001011001000110110;
12'b100111011111: dataA <= 32'b00001101010100110000111101000101;
12'b100111100000: dataA <= 32'b01011001010101100011110111110011;
12'b100111100001: dataA <= 32'b00000010101100010110111000110101;
12'b100111100010: dataA <= 32'b11110110111111001110111000000110;
12'b100111100011: dataA <= 32'b00000000110001010001001010111010;
12'b100111100100: dataA <= 32'b11100000011011000111001000101111;
12'b100111100101: dataA <= 32'b00000111011110001100111010101011;
12'b100111100110: dataA <= 32'b10010110100110111010111001000010;
12'b100111100111: dataA <= 32'b00000100010101001110111101110011;
12'b100111101000: dataA <= 32'b11011011011010000111101000010111;
12'b100111101001: dataA <= 32'b00001001010111011100110001010110;
12'b100111101010: dataA <= 32'b11011111010100101010111000011100;
12'b100111101011: dataA <= 32'b00001101110100110010011000110010;
12'b100111101100: dataA <= 32'b11111100111111011110011100110001;
12'b100111101101: dataA <= 32'b00001001011010010100011110011010;
12'b100111101110: dataA <= 32'b10011001001001101010100101100011;
12'b100111101111: dataA <= 32'b00001000001010100000010001001101;
12'b100111110000: dataA <= 32'b01010101010010101001111111010001;
12'b100111110001: dataA <= 32'b00000110011000001100110001011110;
12'b100111110010: dataA <= 32'b01001001000010001110011000010100;
12'b100111110011: dataA <= 32'b00001100010011100100100000100110;
12'b100111110100: dataA <= 32'b10110010101010001001001010100001;
12'b100111110101: dataA <= 32'b00000101011100010100111110110001;
12'b100111110110: dataA <= 32'b11101101011011110101001011101001;
12'b100111110111: dataA <= 32'b00000111010011011000111001011000;
12'b100111111000: dataA <= 32'b00010011000010111101101000000011;
12'b100111111001: dataA <= 32'b00001011010010111101001101111111;
12'b100111111010: dataA <= 32'b11101100110110001011000111100111;
12'b100111111011: dataA <= 32'b00001000000001100110000111000100;
12'b100111111100: dataA <= 32'b10100011010011011101011111010000;
12'b100111111101: dataA <= 32'b00000001001001011111000000101001;
12'b100111111110: dataA <= 32'b01011000011010110011101011001001;
12'b100111111111: dataA <= 32'b00001001000011110110101010110111;
12'b101000000000: dataA <= 32'b01101010010010001001111010000010;
12'b101000000001: dataA <= 32'b00000101111000010010110010000000;
12'b101000000010: dataA <= 32'b00111001001101011100010011000110;
12'b101000000011: dataA <= 32'b00000100101001100011001010100100;
12'b101000000100: dataA <= 32'b00011110000101011111100001101000;
12'b101000000101: dataA <= 32'b00001000010111011111001010010010;
12'b101000000110: dataA <= 32'b11010100010010110101100111000110;
12'b101000000111: dataA <= 32'b00001010010010011110100010011100;
12'b101000001000: dataA <= 32'b10011001000000010010100011001010;
12'b101000001001: dataA <= 32'b00000010111010001011010010000111;
12'b101000001010: dataA <= 32'b11111101000010111011011010100101;
12'b101000001011: dataA <= 32'b00001001100001111101010111010010;
12'b101000001100: dataA <= 32'b10110000010010011010101101110010;
12'b101000001101: dataA <= 32'b00000110111100001110101010110010;
12'b101000001110: dataA <= 32'b01011011000100001100000010010010;
12'b101000001111: dataA <= 32'b00001010011000100101001101111101;
12'b101000010000: dataA <= 32'b11001110111100101011100110111011;
12'b101000010001: dataA <= 32'b00001110110011110100111000011001;
12'b101000010010: dataA <= 32'b00000000000001010001100111001010;
12'b101000010011: dataA <= 32'b00000000000000000000000000000000;
12'b101000010100: dataA <= 32'b10010100010000010010010010100100;
12'b101000010101: dataA <= 32'b00001000010110011010100110010111;
12'b101000010110: dataA <= 32'b01110010010001000110110011110110;
12'b101000010111: dataA <= 32'b00001101111010111001001110101001;
12'b101000011000: dataA <= 32'b11000010111011000100101100001101;
12'b101000011001: dataA <= 32'b00001011011101101001010000001100;
12'b101000011010: dataA <= 32'b10010110101000101100000101001110;
12'b101000011011: dataA <= 32'b00001010101100101010011001110111;
12'b101000011100: dataA <= 32'b00101000000110100101011010010000;
12'b101000011101: dataA <= 32'b00000100001011001110001111000110;
12'b101000011110: dataA <= 32'b00011010111110000111100111010111;
12'b101000011111: dataA <= 32'b00001001110110011110000101101101;
12'b101000100000: dataA <= 32'b10100100110111000011111101101010;
12'b101000100001: dataA <= 32'b00001000100110110001011010010100;
12'b101000100010: dataA <= 32'b01010001100111010011001101000110;
12'b101000100011: dataA <= 32'b00001100111011101000101100001101;
12'b101000100100: dataA <= 32'b00011011100001011110010111010011;
12'b101000100101: dataA <= 32'b00000101000001100101011000100011;
12'b101000100110: dataA <= 32'b00111010111111101101111101000101;
12'b101000100111: dataA <= 32'b00001010110101110101101111100101;
12'b101000101000: dataA <= 32'b10010100011111000100101111010000;
12'b101000101001: dataA <= 32'b00001010110011101000011100100001;
12'b101000101010: dataA <= 32'b11010100111001111011111001010101;
12'b101000101011: dataA <= 32'b00001011111100100000001001011100;
12'b101000101100: dataA <= 32'b11100100000101000111010110111110;
12'b101000101101: dataA <= 32'b00001010010010101101011110111100;
12'b101000101110: dataA <= 32'b01001100101010000010011010010101;
12'b101000101111: dataA <= 32'b00001010000001110100010100001011;
12'b101000110000: dataA <= 32'b00010011001010001110000110100011;
12'b101000110001: dataA <= 32'b00001000111110011100111100110011;
12'b101000110010: dataA <= 32'b11000010111101011111100101111000;
12'b101000110011: dataA <= 32'b00000110011100010111010000101110;
12'b101000110100: dataA <= 32'b01001000010100010010010111110110;
12'b101000110101: dataA <= 32'b00001100110110110001000100111101;
12'b101000110110: dataA <= 32'b11010111010001100011100111010011;
12'b101000110111: dataA <= 32'b00000011001010011000111000101100;
12'b101000111000: dataA <= 32'b01110111000110111111011001000110;
12'b101000111001: dataA <= 32'b00000000101110010001000111000011;
12'b101000111010: dataA <= 32'b00100100011010110111011000101111;
12'b101000111011: dataA <= 32'b00000101111110001110110010101100;
12'b101000111100: dataA <= 32'b10011000100011000011011010100010;
12'b101000111101: dataA <= 32'b00000011110011010000111001110011;
12'b101000111110: dataA <= 32'b10011001011001101111100111110111;
12'b101000111111: dataA <= 32'b00001000011000011100110001000110;
12'b101001000000: dataA <= 32'b10011101010100110010010111011011;
12'b101001000001: dataA <= 32'b00001101010110110110100000111010;
12'b101001000010: dataA <= 32'b00111101000111001110111100010011;
12'b101001000011: dataA <= 32'b00001000011010011000011010100011;
12'b101001000100: dataA <= 32'b01011001001001110010100111000010;
12'b101001000101: dataA <= 32'b00001000101010100100010001000101;
12'b101001000110: dataA <= 32'b00010011001010111010001111010100;
12'b101001000111: dataA <= 32'b00000101110111001100101001010110;
12'b101001001000: dataA <= 32'b11001000111001111110010111110100;
12'b101001001001: dataA <= 32'b00001011110100101000100100010101;
12'b101001001010: dataA <= 32'b00110100110010100001011011100011;
12'b101001001011: dataA <= 32'b00000011111010010100111011000010;
12'b101001001100: dataA <= 32'b10101011011111100101111100001011;
12'b101001001101: dataA <= 32'b00000110110010011010110101110000;
12'b101001001110: dataA <= 32'b00010010111010110101111001000011;
12'b101001001111: dataA <= 32'b00001011010011111011010101101111;
12'b101001010000: dataA <= 32'b00101100111010010011011000100111;
12'b101001010001: dataA <= 32'b00001001100001101100001010111101;
12'b101001010010: dataA <= 32'b01100001010111010101111111010010;
12'b101001010011: dataA <= 32'b00000001100111011111000000111001;
12'b101001010100: dataA <= 32'b10011100011010110100001011101010;
12'b101001010101: dataA <= 32'b00001010000100111000110110011111;
12'b101001010110: dataA <= 32'b01101110010110010001111011000011;
12'b101001010111: dataA <= 32'b00000100110111010100101110011000;
12'b101001011000: dataA <= 32'b01110111010101010100000100000100;
12'b101001011001: dataA <= 32'b00000101001000100001001010100100;
12'b101001011010: dataA <= 32'b01100100000101000111010010000110;
12'b101001011011: dataA <= 32'b00000111110111011101001010100010;
12'b101001011100: dataA <= 32'b00011010001110101101111000000110;
12'b101001011101: dataA <= 32'b00001010010010100000100010010101;
12'b101001011110: dataA <= 32'b10011000111100011001110011101001;
12'b101001011111: dataA <= 32'b00000001110111001011001001101111;
12'b101001100000: dataA <= 32'b01111101001010111011101011100111;
12'b101001100001: dataA <= 32'b00001010100010111001011111010011;
12'b101001100010: dataA <= 32'b11110100011010100010111101010101;
12'b101001100011: dataA <= 32'b00000101111011010000100010111010;
12'b101001100100: dataA <= 32'b01011011000000001011010010010000;
12'b101001100101: dataA <= 32'b00001001011001100101001101110101;
12'b101001100110: dataA <= 32'b01010000111000101011000101011010;
12'b101001100111: dataA <= 32'b00001110010101110101000000101001;
12'b101001101000: dataA <= 32'b00000000000001100001010111101001;
12'b101001101001: dataA <= 32'b00000000000000000000000000000000;
12'b101001101010: dataA <= 32'b10011000001100011001110100000011;
12'b101001101011: dataA <= 32'b00000111110110011100100101111111;
12'b101001101100: dataA <= 32'b10110110011000101110100011010100;
12'b101001101101: dataA <= 32'b00001100011100110111010110111001;
12'b101001101110: dataA <= 32'b00000010101110111101001100001111;
12'b101001101111: dataA <= 32'b00001001111110100111010100001100;
12'b101001110000: dataA <= 32'b10011000100100101011010101001101;
12'b101001110001: dataA <= 32'b00001010101101101110100001011111;
12'b101001110010: dataA <= 32'b10101110001010011101101010010001;
12'b101001110011: dataA <= 32'b00000100101001010010001010111110;
12'b101001110100: dataA <= 32'b00011010111101101111100110010111;
12'b101001110101: dataA <= 32'b00001001010110100100000101100101;
12'b101001110110: dataA <= 32'b10100100110111000100011110001100;
12'b101001110111: dataA <= 32'b00001001100110101101100010010100;
12'b101001111000: dataA <= 32'b10001101011111010011101110001000;
12'b101001111001: dataA <= 32'b00001011011101101010110000001100;
12'b101001111010: dataA <= 32'b10010111011101001110000110110011;
12'b101001111011: dataA <= 32'b00000110100001100011011000101010;
12'b101001111100: dataA <= 32'b10111011000111011110011110000111;
12'b101001111101: dataA <= 32'b00001010010110101111110011011101;
12'b101001111110: dataA <= 32'b00011000011010111101001111010011;
12'b101001111111: dataA <= 32'b00001010010100101100100000110001;
12'b101010000000: dataA <= 32'b10010100110101111011111000110101;
12'b101010000001: dataA <= 32'b00001010111110100100001001011100;
12'b101010000010: dataA <= 32'b00101010001000110110110101111110;
12'b101010000011: dataA <= 32'b00001001110011101001100010110101;
12'b101010000100: dataA <= 32'b11010000100010001010011001110110;
12'b101010000101: dataA <= 32'b00001011100011111000011100001010;
12'b101010000110: dataA <= 32'b10010011000101111110010111100010;
12'b101010000111: dataA <= 32'b00000111011110011100111100111010;
12'b101010001000: dataA <= 32'b00000010110001000111010100110111;
12'b101010001001: dataA <= 32'b00000101011011010101001100011110;
12'b101010001010: dataA <= 32'b11001110001100011001110111010110;
12'b101010001011: dataA <= 32'b00001011111000110001001100110100;
12'b101010001100: dataA <= 32'b01010101001101100011100111010011;
12'b101010001101: dataA <= 32'b00000011101000011000110100101100;
12'b101010001110: dataA <= 32'b11110101001110100111101010000111;
12'b101010001111: dataA <= 32'b00000000101011001110111111000011;
12'b101010010000: dataA <= 32'b01101000011110011111101000101111;
12'b101010010001: dataA <= 32'b00000100011101010000101010101100;
12'b101010010010: dataA <= 32'b10011100100011000011111011100100;
12'b101010010011: dataA <= 32'b00000011110001010000110001110011;
12'b101010010100: dataA <= 32'b00010111010101011111100110110111;
12'b101010010101: dataA <= 32'b00000111011000011110110000110110;
12'b101010010110: dataA <= 32'b00011011010101000001110110011011;
12'b101010010111: dataA <= 32'b00001100011000111000101001001010;
12'b101010011000: dataA <= 32'b01111011010010110111011011110101;
12'b101010011001: dataA <= 32'b00000110111010011100011010100011;
12'b101010011010: dataA <= 32'b11011001000101111010101000000010;
12'b101010011011: dataA <= 32'b00001001001010101000010100111100;
12'b101010011100: dataA <= 32'b10010011000111000010101110110111;
12'b101010011101: dataA <= 32'b00000100110110010000100001000101;
12'b101010011110: dataA <= 32'b00001010110001101110010111010100;
12'b101010011111: dataA <= 32'b00001011010110101010101000001101;
12'b101010100000: dataA <= 32'b10110100111010110001101101000101;
12'b101010100001: dataA <= 32'b00000010111001010100110111001010;
12'b101010100010: dataA <= 32'b10100111100011011110011100101101;
12'b101010100011: dataA <= 32'b00000110110010011010110110000000;
12'b101010100100: dataA <= 32'b11010010110110100110001010000100;
12'b101010100101: dataA <= 32'b00001010110100111001100001011110;
12'b101010100110: dataA <= 32'b10101111000010010011011001100111;
12'b101010100111: dataA <= 32'b00001011000010110000001110110101;
12'b101010101000: dataA <= 32'b11011111010111000110011110110101;
12'b101010101001: dataA <= 32'b00000010100101011111000001001000;
12'b101010101010: dataA <= 32'b10100000010110110100011100001100;
12'b101010101011: dataA <= 32'b00001011000101111010111110000111;
12'b101010101100: dataA <= 32'b10110010011110100010001100000101;
12'b101010101101: dataA <= 32'b00000100010101010110101010110000;
12'b101010101110: dataA <= 32'b10110011100001010011110101000011;
12'b101010101111: dataA <= 32'b00000110000111100001001010100100;
12'b101010110000: dataA <= 32'b10101010001000110110110011000100;
12'b101010110001: dataA <= 32'b00000110110111011101001010101010;
12'b101010110010: dataA <= 32'b00011110001010011110001001000110;
12'b101010110011: dataA <= 32'b00001001110011100100100010001101;
12'b101010110100: dataA <= 32'b10011000111100101001010100100111;
12'b101010110101: dataA <= 32'b00000000110101001001000001011111;
12'b101010110110: dataA <= 32'b11111011010111000100001100101001;
12'b101010110111: dataA <= 32'b00001100000011110101101011011011;
12'b101010111000: dataA <= 32'b01111000100010101011001100110111;
12'b101010111001: dataA <= 32'b00000100111010010100011110111011;
12'b101010111010: dataA <= 32'b01011011000000010010100010001110;
12'b101010111011: dataA <= 32'b00001000011001100011001101101101;
12'b101010111100: dataA <= 32'b11010000110000110010100100011001;
12'b101010111101: dataA <= 32'b00001101010111110101001100111000;
12'b101010111110: dataA <= 32'b00000000000001110001011000001001;
12'b101010111111: dataA <= 32'b00000000000000000000000000000000;
endcase
if (enB)
case(addrB)
12'b000000000000: dataB <= 32'b00000111001100111111000001110111;
12'b000000000001: dataB <= 32'b00001011010000010011000111110100;
12'b000000000010: dataB <= 32'b00001100010011010110101010011001;
12'b000000000011: dataB <= 32'b00001110000111101010010000110010;
12'b000000000100: dataB <= 32'b10010111111010100010000111100111;
12'b000000000101: dataB <= 32'b00001111001100101010110010000111;
12'b000000000110: dataB <= 32'b00010011001101101110100110110101;
12'b000000000111: dataB <= 32'b00000110101010010000100011110101;
12'b000000001000: dataB <= 32'b00000100100010110011001000101011;
12'b000000001001: dataB <= 32'b00000100110110000101011011010010;
12'b000000001010: dataB <= 32'b11011111001011110100101011110011;
12'b000000001011: dataB <= 32'b00001011001101000010110110100100;
12'b000000001100: dataB <= 32'b01011010110110001001110110000011;
12'b000000001101: dataB <= 32'b00000011001100110000100110010011;
12'b000000001110: dataB <= 32'b10101111100101110001010100000011;
12'b000000001111: dataB <= 32'b00001110101001011000101010010111;
12'b000000010000: dataB <= 32'b10101111010011000101101001110010;
12'b000000010001: dataB <= 32'b00000000110010101100111001010110;
12'b000000010010: dataB <= 32'b00100010001011001001000011100011;
12'b000000010011: dataB <= 32'b00001011001011111000100010110001;
12'b000000010100: dataB <= 32'b01001101001110100010001001100001;
12'b000000010101: dataB <= 32'b00001010001011010000100100100110;
12'b000000010110: dataB <= 32'b00011011010101111100001010101110;
12'b000000010111: dataB <= 32'b00001111001010000100110110010101;
12'b000000011000: dataB <= 32'b01000100101011011110011111010100;
12'b000000011001: dataB <= 32'b00001001101100110000101110100010;
12'b000000011010: dataB <= 32'b10010001011101001011101011001100;
12'b000000011011: dataB <= 32'b00000001101000001110001101011111;
12'b000000011100: dataB <= 32'b00100011011011001100000001010000;
12'b000000011101: dataB <= 32'b00001111010001011111000101010110;
12'b000000011110: dataB <= 32'b00011001111011101101111011110110;
12'b000000011111: dataB <= 32'b00001101110101100111010111000111;
12'b000000100000: dataB <= 32'b01000111100000111111001011010001;
12'b000000100001: dataB <= 32'b00001100001000100110011110011110;
12'b000000100010: dataB <= 32'b10100111010101110100111001110001;
12'b000000100011: dataB <= 32'b00000100011000011011001110001110;
12'b000000100100: dataB <= 32'b11100110010111110010110011101011;
12'b000000100101: dataB <= 32'b00000101111110011111100001111001;
12'b000000100110: dataB <= 32'b10001110101111110011000111101110;
12'b000000100111: dataB <= 32'b00001110110111010101011110001010;
12'b000000101000: dataB <= 32'b01010001000101111001110010001000;
12'b000000101001: dataB <= 32'b00001000111000011001011101110100;
12'b000000101010: dataB <= 32'b01101011010011110101001011110010;
12'b000000101011: dataB <= 32'b00001100010001011001000011000110;
12'b000000101100: dataB <= 32'b10101011001000111101111101110011;
12'b000000101101: dataB <= 32'b00001100000111010100001101000101;
12'b000000101110: dataB <= 32'b11101000001011101010011010101000;
12'b000000101111: dataB <= 32'b00001101010010001101000101101010;
12'b000000110000: dataB <= 32'b00100011001101010100000001001111;
12'b000000110001: dataB <= 32'b00000101001101001010101110011110;
12'b000000110010: dataB <= 32'b11100011011001010001111011100010;
12'b000000110011: dataB <= 32'b00001011010110010001011110110101;
12'b000000110100: dataB <= 32'b10011001101011001100101010010001;
12'b000000110101: dataB <= 32'b00001011001001010100101010100111;
12'b000000110110: dataB <= 32'b10011100010100110010010010100101;
12'b000000110111: dataB <= 32'b00001100111010011011010101010001;
12'b000000111000: dataB <= 32'b11110000110011001001000110100110;
12'b000000111001: dataB <= 32'b00001001010010011011001000010011;
12'b000000111010: dataB <= 32'b00011011011011000010110010001011;
12'b000000111011: dataB <= 32'b00001010001010110000001111011101;
12'b000000111100: dataB <= 32'b01100000100001101011010011101100;
12'b000000111101: dataB <= 32'b00000001001001000110011110110010;
12'b000000111110: dataB <= 32'b10101011000011001001111010100010;
12'b000000111111: dataB <= 32'b00000010111010100001000000011101;
12'b000001000000: dataB <= 32'b11001010111110001010010110000111;
12'b000001000001: dataB <= 32'b00000010101001011110001011110011;
12'b000001000010: dataB <= 32'b01001110011001000010110010100111;
12'b000001000011: dataB <= 32'b00001010110111010101010000010010;
12'b000001000100: dataB <= 32'b11110000011001111101010001110101;
12'b000001000101: dataB <= 32'b00000011110011100100111110010010;
12'b000001000110: dataB <= 32'b10000100101011011110010010011001;
12'b000001000111: dataB <= 32'b00001011110010100101000101010010;
12'b000001001000: dataB <= 32'b10000101000011000011000011001101;
12'b000001001001: dataB <= 32'b00001001101100010000110110100011;
12'b000001001010: dataB <= 32'b00011111001100101110100011110110;
12'b000001001011: dataB <= 32'b00001010111110100001101111110101;
12'b000001001100: dataB <= 32'b00101010001010000001110100100110;
12'b000001001101: dataB <= 32'b00000001100111110100010101111001;
12'b000001001110: dataB <= 32'b00010000001101100010101011100110;
12'b000001001111: dataB <= 32'b00001101010110001111010101101010;
12'b000001010000: dataB <= 32'b10100001001001010111010111011011;
12'b000001010001: dataB <= 32'b00001100101111100110111010101100;
12'b000001010010: dataB <= 32'b00011001011101010110011100110111;
12'b000001010011: dataB <= 32'b00001011100101100110010100011110;
12'b000001010100: dataB <= 32'b00000000000000101100010100101111;
12'b000001010101: dataB <= 32'b00000000000000000000000000000000;
12'b000001010110: dataB <= 32'b01001001010101001111010010011010;
12'b000001010111: dataB <= 32'b00001011001111010011001011110011;
12'b000001011000: dataB <= 32'b10001000011011011101111011011000;
12'b000001011001: dataB <= 32'b00001101000100100110001100101010;
12'b000001011010: dataB <= 32'b10011101111010010001110110100111;
12'b000001011011: dataB <= 32'b00001110101001101000101110011111;
12'b000001011100: dataB <= 32'b01010101010010000110100111010101;
12'b000001011101: dataB <= 32'b00000110001010001100101011110100;
12'b000001011110: dataB <= 32'b11000010101110101010111000001011;
12'b000001011111: dataB <= 32'b00000101110111000111100011000001;
12'b000001100000: dataB <= 32'b10011111001011110011111011110001;
12'b000001100001: dataB <= 32'b00001011001100000011000010100100;
12'b000001100010: dataB <= 32'b01011010110101111001110101000100;
12'b000001100011: dataB <= 32'b00000011001110101100011110010011;
12'b000001100100: dataB <= 32'b10110011011101100001010011000101;
12'b000001100101: dataB <= 32'b00001101100110010110101110101111;
12'b000001100110: dataB <= 32'b11110001001011001101001001110001;
12'b000001100111: dataB <= 32'b00000000110101101100110101100110;
12'b000001101000: dataB <= 32'b11011110001010111000100010100101;
12'b000001101001: dataB <= 32'b00001010101010110110010110100000;
12'b000001101010: dataB <= 32'b11001111010110010001111000000001;
12'b000001101011: dataB <= 32'b00001001101010001110101100110110;
12'b000001101100: dataB <= 32'b00011101010101111100001010101101;
12'b000001101101: dataB <= 32'b00001110001000000100111110011101;
12'b000001101110: dataB <= 32'b00000010110111101101111111010010;
12'b000001101111: dataB <= 32'b00001001001011101110100110011010;
12'b000001110000: dataB <= 32'b10010101100101001011111010101011;
12'b000001110001: dataB <= 32'b00000000101011001010010101101111;
12'b000001110010: dataB <= 32'b01100101011011000011100001110010;
12'b000001110011: dataB <= 32'b00001111001110011111000101100110;
12'b000001110100: dataB <= 32'b10011111111011110101001100010100;
12'b000001110101: dataB <= 32'b00001110010011101001010011011110;
12'b000001110110: dataB <= 32'b00001011101101001111011011010000;
12'b000001110111: dataB <= 32'b00001011000110100010011110101110;
12'b000001111000: dataB <= 32'b10101001010001110100111001110001;
12'b000001111001: dataB <= 32'b00000101011001011101001110011110;
12'b000001111010: dataB <= 32'b11100010010011101010000011001101;
12'b000001111011: dataB <= 32'b00000111011110100011011101101001;
12'b000001111100: dataB <= 32'b10001100110111101010010111101110;
12'b000001111101: dataB <= 32'b00001111010100011001100010000010;
12'b000001111110: dataB <= 32'b01010001001101101001110001001010;
12'b000001111111: dataB <= 32'b00001001111000011101011101110100;
12'b000010000000: dataB <= 32'b11101101001111110100101011110000;
12'b000010000001: dataB <= 32'b00001100001111011001000111010101;
12'b000010000010: dataB <= 32'b00101011000101001110011101110001;
12'b000010000011: dataB <= 32'b00001011000101010000010001010110;
12'b000010000100: dataB <= 32'b11100010000111011001101001100111;
12'b000010000101: dataB <= 32'b00001101001111001101001101100010;
12'b000010000110: dataB <= 32'b11100101001101010100010001010001;
12'b000010000111: dataB <= 32'b00000101001110001000110110101101;
12'b000010001000: dataB <= 32'b01100101011001000010001010000001;
12'b000010001001: dataB <= 32'b00001011110100010101100111000101;
12'b000010001010: dataB <= 32'b01011101101111001100001010010000;
12'b000010001011: dataB <= 32'b00001010001000010010101110111111;
12'b000010001100: dataB <= 32'b11011000010100101010110001101000;
12'b000010001101: dataB <= 32'b00001101011000011101010101000001;
12'b000010001110: dataB <= 32'b01101110101010111000110101100111;
12'b000010001111: dataB <= 32'b00001001010010011011001000010100;
12'b000010010000: dataB <= 32'b10011101011010111010010001101101;
12'b000010010001: dataB <= 32'b00001001101001101010001011100100;
12'b000010010010: dataB <= 32'b00011100100101101011010011101110;
12'b000010010011: dataB <= 32'b00000000101100000100100110100010;
12'b000010010100: dataB <= 32'b00101010111110111001011001000001;
12'b000010010101: dataB <= 32'b00000011111100100001000000101110;
12'b000010010110: dataB <= 32'b00001101000110000010010101001000;
12'b000010010111: dataB <= 32'b00000010001011011010001111110011;
12'b000010011000: dataB <= 32'b00001010100000111011010001101001;
12'b000010011001: dataB <= 32'b00001011110110010111010100001011;
12'b000010011010: dataB <= 32'b11101010010010000101010010010111;
12'b000010011011: dataB <= 32'b00000100010101100100111110001010;
12'b000010011100: dataB <= 32'b11000010110111101101110011011011;
12'b000010011101: dataB <= 32'b00001011110000100101000101001010;
12'b000010011110: dataB <= 32'b01000111001010111010100011001111;
12'b000010011111: dataB <= 32'b00001001001011010000111110100011;
12'b000010100000: dataB <= 32'b10011111001100111111000100111000;
12'b000010100001: dataB <= 32'b00001011111100100101101011110100;
12'b000010100010: dataB <= 32'b01100100000101110010000011101000;
12'b000010100011: dataB <= 32'b00000001001010101110001101101001;
12'b000010100100: dataB <= 32'b00001100010101011010111010100101;
12'b000010100101: dataB <= 32'b00001101110100010001011101011010;
12'b000010100110: dataB <= 32'b01100001001001101111101000011011;
12'b000010100111: dataB <= 32'b00001100101101100110110110101100;
12'b000010101000: dataB <= 32'b10011101011101100110101101010101;
12'b000010101001: dataB <= 32'b00001010100011100000010100101110;
12'b000010101010: dataB <= 32'b00000000000000101100110100110000;
12'b000010101011: dataB <= 32'b00000000000000000000000000000000;
12'b000010101100: dataB <= 32'b10001011011101100111100011111100;
12'b000010101101: dataB <= 32'b00001010101110010101010011110010;
12'b000010101110: dataB <= 32'b01000110100011101101011100010110;
12'b000010101111: dataB <= 32'b00001011100011100000001000100011;
12'b000010110000: dataB <= 32'b01100011111010001001110101101000;
12'b000010110001: dataB <= 32'b00001110000111100110101010110111;
12'b000010110010: dataB <= 32'b10010111010110010110100111110101;
12'b000010110011: dataB <= 32'b00000101101011001100110011110011;
12'b000010110100: dataB <= 32'b01000010111010100010100111101011;
12'b000010110101: dataB <= 32'b00000110011000001011101010110001;
12'b000010110110: dataB <= 32'b01100001001011110011001100010000;
12'b000010110111: dataB <= 32'b00001010101010000011001110101100;
12'b000010111000: dataB <= 32'b00011000111001101010000100000101;
12'b000010111001: dataB <= 32'b00000011010000101010011010001011;
12'b000010111010: dataB <= 32'b00110101010101010001100010000111;
12'b000010111011: dataB <= 32'b00001100100100010100110010111111;
12'b000010111100: dataB <= 32'b00110001000111010100101010010001;
12'b000010111101: dataB <= 32'b00000001110111101010101101110111;
12'b000010111110: dataB <= 32'b10011000001110100000010001100111;
12'b000010111111: dataB <= 32'b00001010001001110000001110001000;
12'b000011000000: dataB <= 32'b00010001011110001001110110100001;
12'b000011000001: dataB <= 32'b00001001001010001100110101000111;
12'b000011000010: dataB <= 32'b11011111010101111100001010001100;
12'b000011000011: dataB <= 32'b00001101000101000101001010100100;
12'b000011000100: dataB <= 32'b00000010111111110101001111001111;
12'b000011000101: dataB <= 32'b00001001001011101100100010001010;
12'b000011000110: dataB <= 32'b10011001100101001100011010001010;
12'b000011000111: dataB <= 32'b00000000101101000110011110000111;
12'b000011001000: dataB <= 32'b01101001010111000011000010010101;
12'b000011001001: dataB <= 32'b00001111001011011111000101110110;
12'b000011001010: dataB <= 32'b11100101111011110100011100110010;
12'b000011001011: dataB <= 32'b00001110110000101011001111100101;
12'b000011001100: dataB <= 32'b11010001110001100111101011001110;
12'b000011001101: dataB <= 32'b00001010000101011110011110111101;
12'b000011001110: dataB <= 32'b01101011001101111100111001110000;
12'b000011001111: dataB <= 32'b00000110011010011101010010101110;
12'b000011010000: dataB <= 32'b00011110010011011001100011001111;
12'b000011010001: dataB <= 32'b00001000111110100101011101011010;
12'b000011010010: dataB <= 32'b10001100111111100001110111101110;
12'b000011010011: dataB <= 32'b00001111010001011101100101111010;
12'b000011010100: dataB <= 32'b01010011010001011010000001001101;
12'b000011010101: dataB <= 32'b00001010110111011111100001110100;
12'b000011010110: dataB <= 32'b01101101001011110011111011101111;
12'b000011010111: dataB <= 32'b00001011101101011001000111011101;
12'b000011011000: dataB <= 32'b01101011000001011110101110001111;
12'b000011011001: dataB <= 32'b00001010000100001100011001011110;
12'b000011011010: dataB <= 32'b00011110000111001001001000100110;
12'b000011011011: dataB <= 32'b00001101001101001111010101011011;
12'b000011011100: dataB <= 32'b10100101001101010100100001110100;
12'b000011011101: dataB <= 32'b00000101001111001000111110110101;
12'b000011011110: dataB <= 32'b00101001010100111010101000100001;
12'b000011011111: dataB <= 32'b00001100010011011001100111001101;
12'b000011100000: dataB <= 32'b11100001101111001011101010001111;
12'b000011100001: dataB <= 32'b00001001100111010000110111001110;
12'b000011100010: dataB <= 32'b01010100011000100011100000101010;
12'b000011100011: dataB <= 32'b00001110010101011111010100110010;
12'b000011100100: dataB <= 32'b00101100100110100000010100101000;
12'b000011100101: dataB <= 32'b00001001110001011101001100011101;
12'b000011100110: dataB <= 32'b00100001011010110010000001101111;
12'b000011100111: dataB <= 32'b00001001001001100110000111100100;
12'b000011101000: dataB <= 32'b11011010100101100011100011110000;
12'b000011101001: dataB <= 32'b00000000101111000010110010011001;
12'b000011101010: dataB <= 32'b10101000111010101001001000000001;
12'b000011101011: dataB <= 32'b00000100111101100001000000110110;
12'b000011101100: dataB <= 32'b01001101001101110010010100101001;
12'b000011101101: dataB <= 32'b00000001101101010100010011101010;
12'b000011101110: dataB <= 32'b11001000101000111011100001001011;
12'b000011101111: dataB <= 32'b00001100010100011001011000001011;
12'b000011110000: dataB <= 32'b11100110001110001101000011011001;
12'b000011110001: dataB <= 32'b00000100110110100100111010000010;
12'b000011110010: dataB <= 32'b01000011000011110101000100011100;
12'b000011110011: dataB <= 32'b00001011101111100101000001000011;
12'b000011110100: dataB <= 32'b00001001010110110010010011010001;
12'b000011110101: dataB <= 32'b00001001001011010001000010011011;
12'b000011110110: dataB <= 32'b11100001001101010111010101011001;
12'b000011110111: dataB <= 32'b00001101011010101001101011110011;
12'b000011111000: dataB <= 32'b01100000000101101010000010101010;
12'b000011111001: dataB <= 32'b00000000101100101010000101011001;
12'b000011111010: dataB <= 32'b01001000011101010011001001000100;
12'b000011111011: dataB <= 32'b00001110010010010101100001010010;
12'b000011111100: dataB <= 32'b00100011001010000111101001011011;
12'b000011111101: dataB <= 32'b00001100001011100110110110101100;
12'b000011111110: dataB <= 32'b00011111100001110110101101110010;
12'b000011111111: dataB <= 32'b00001001100010011100010100111111;
12'b000100000000: dataB <= 32'b00000000000000110101010101010001;
12'b000100000001: dataB <= 32'b00000000000000000000000000000000;
12'b000100000010: dataB <= 32'b00001111100101111111100100111101;
12'b000100000011: dataB <= 32'b00001010101100010111010111100010;
12'b000100000100: dataB <= 32'b11000010101111101100101100110101;
12'b000100000101: dataB <= 32'b00001010100001011100001100011011;
12'b000100000110: dataB <= 32'b00101001111001111001110101001001;
12'b000100000111: dataB <= 32'b00001101000101100100100111000111;
12'b000100001000: dataB <= 32'b11011001011010100110011000010101;
12'b000100001001: dataB <= 32'b00000101001100001010111011110010;
12'b000100001010: dataB <= 32'b00000011000110011010010111101011;
12'b000100001011: dataB <= 32'b00000111011001010001110010100001;
12'b000100001100: dataB <= 32'b00100001001011101010011011101110;
12'b000100001101: dataB <= 32'b00001010001010000101011010101100;
12'b000100001110: dataB <= 32'b00011000111001100010000011000111;
12'b000100001111: dataB <= 32'b00000011010010100110010110001011;
12'b000100010000: dataB <= 32'b10110111001101001001110001101001;
12'b000100010001: dataB <= 32'b00001011100010010010110111010110;
12'b000100010010: dataB <= 32'b00110000111111010100001010010000;
12'b000100010011: dataB <= 32'b00000010111010101000101010000111;
12'b000100010100: dataB <= 32'b10010100010010001000010001001010;
12'b000100010101: dataB <= 32'b00001001001000101100001001111000;
12'b000100010110: dataB <= 32'b10010101100001111001110101000001;
12'b000100010111: dataB <= 32'b00001000101001001100111101011111;
12'b000100011000: dataB <= 32'b10100001010101111100001010001011;
12'b000100011001: dataB <= 32'b00001100000011000111010110100100;
12'b000100011010: dataB <= 32'b00000011001011110100011111001100;
12'b000100011011: dataB <= 32'b00001000101011101000011110000010;
12'b000100011100: dataB <= 32'b10011101101001010100101001101001;
12'b000100011101: dataB <= 32'b00000000110000000100101010011111;
12'b000100011110: dataB <= 32'b01101011010010111010110010110111;
12'b000100011111: dataB <= 32'b00001110101000011111000110000110;
12'b000100100000: dataB <= 32'b01101011111011110011101100110000;
12'b000100100001: dataB <= 32'b00001110001110101101001011110101;
12'b000100100010: dataB <= 32'b01010101111001111111101010101101;
12'b000100100011: dataB <= 32'b00001001000100011100011111000101;
12'b000100100100: dataB <= 32'b00101101001010000100111001101111;
12'b000100100101: dataB <= 32'b00000111011011011111010010110110;
12'b000100100110: dataB <= 32'b01011010010111001001000011010001;
12'b000100100111: dataB <= 32'b00001010011110101001011001010010;
12'b000100101000: dataB <= 32'b10001101000111010001010111001110;
12'b000100101001: dataB <= 32'b00001111001110011111100101110010;
12'b000100101010: dataB <= 32'b10010101010101010010010000110000;
12'b000100101011: dataB <= 32'b00001011010110100011011101111100;
12'b000100101100: dataB <= 32'b10101111000011110011001011101101;
12'b000100101101: dataB <= 32'b00001011101100011001001011100100;
12'b000100101110: dataB <= 32'b01101010111101101110111101101100;
12'b000100101111: dataB <= 32'b00001000100100001000100001101110;
12'b000100110000: dataB <= 32'b01011000001010111000101000000110;
12'b000100110001: dataB <= 32'b00001100101011010001011101011011;
12'b000100110010: dataB <= 32'b01100111001001011100110010010110;
12'b000100110011: dataB <= 32'b00000101010000001001000111000101;
12'b000100110100: dataB <= 32'b10101011010000110011000111000001;
12'b000100110101: dataB <= 32'b00001100110001011101101011001100;
12'b000100110110: dataB <= 32'b01100101101011000011001010001111;
12'b000100110111: dataB <= 32'b00001000100110010000111011011110;
12'b000100111000: dataB <= 32'b11010010011100100100000000101101;
12'b000100111001: dataB <= 32'b00001110110011100001010100101010;
12'b000100111010: dataB <= 32'b10101010011110010000010100001001;
12'b000100111011: dataB <= 32'b00001001110001011101001100100101;
12'b000100111100: dataB <= 32'b01100011011010100001110001110010;
12'b000100111101: dataB <= 32'b00001000001000100000000111100011;
12'b000100111110: dataB <= 32'b10011000100101100011100011110001;
12'b000100111111: dataB <= 32'b00000000110010000010111110001001;
12'b000101000000: dataB <= 32'b00101000110110010000110110100001;
12'b000101000001: dataB <= 32'b00000110011110100001000001001111;
12'b000101000010: dataB <= 32'b11001111010101101010100011101010;
12'b000101000011: dataB <= 32'b00000001110000010000010111100001;
12'b000101000100: dataB <= 32'b10000110110100111100000000101110;
12'b000101000101: dataB <= 32'b00001100010011011011011000001100;
12'b000101000110: dataB <= 32'b11100010001110010101000100011011;
12'b000101000111: dataB <= 32'b00000101011000100100111001111010;
12'b000101001000: dataB <= 32'b10000011001011110100010101111110;
12'b000101001001: dataB <= 32'b00001011101101100101000001000011;
12'b000101001010: dataB <= 32'b00001011011110101001110011110011;
12'b000101001011: dataB <= 32'b00001000101011010001001010011011;
12'b000101001100: dataB <= 32'b00100011001001101111100110011010;
12'b000101001101: dataB <= 32'b00001110011000101101100111110011;
12'b000101001110: dataB <= 32'b10011010000101011010010010101100;
12'b000101001111: dataB <= 32'b00000000101111100100000101001001;
12'b000101010000: dataB <= 32'b11000110100101001011011000000011;
12'b000101010001: dataB <= 32'b00001110001111011001100101001010;
12'b000101010010: dataB <= 32'b11100011001010010111101010011010;
12'b000101010011: dataB <= 32'b00001011101001100100110010101011;
12'b000101010100: dataB <= 32'b01100011011110001110101110010000;
12'b000101010101: dataB <= 32'b00001000000010011000010101010111;
12'b000101010110: dataB <= 32'b00000000000000111101100101010011;
12'b000101010111: dataB <= 32'b00000000000000000000000000000000;
12'b000101011000: dataB <= 32'b01010011101110010111100110011110;
12'b000101011001: dataB <= 32'b00001010001011011001011011010001;
12'b000101011010: dataB <= 32'b01000010110111110100001101010011;
12'b000101011011: dataB <= 32'b00001001000001010110001100100100;
12'b000101011100: dataB <= 32'b10101111110101101001110100101010;
12'b000101011101: dataB <= 32'b00001011100011100010100111010110;
12'b000101011110: dataB <= 32'b00011011011110101110001000110101;
12'b000101011111: dataB <= 32'b00000101001101001011000011101010;
12'b000101100000: dataB <= 32'b11000011010010010010000111001011;
12'b000101100001: dataB <= 32'b00001000011001010101111010010000;
12'b000101100010: dataB <= 32'b11100001001011100001111011101101;
12'b000101100011: dataB <= 32'b00001001001001000111100010101011;
12'b000101100100: dataB <= 32'b00011000111101011010010010001001;
12'b000101100101: dataB <= 32'b00000011110100100010010110000011;
12'b000101100110: dataB <= 32'b00111001000000111010010001001100;
12'b000101100111: dataB <= 32'b00001010000001010010111011100110;
12'b000101101000: dataB <= 32'b11110000110111010011101010001111;
12'b000101101001: dataB <= 32'b00000011111100100110100110011110;
12'b000101101010: dataB <= 32'b10001110010101110000010000101101;
12'b000101101011: dataB <= 32'b00001000101000100110000101100000;
12'b000101101100: dataB <= 32'b10010111100101101001110100000011;
12'b000101101101: dataB <= 32'b00001000001001001101000001101111;
12'b000101101110: dataB <= 32'b01100011010101111100001001101010;
12'b000101101111: dataB <= 32'b00001011000010001001011110101100;
12'b000101110000: dataB <= 32'b00000101010111110011101110101001;
12'b000101110001: dataB <= 32'b00001000001011100100011001110010;
12'b000101110010: dataB <= 32'b01100001101001010100111001001000;
12'b000101110011: dataB <= 32'b00000000110011000010110110110111;
12'b000101110100: dataB <= 32'b01101101001110110010010011011001;
12'b000101110101: dataB <= 32'b00001101100110100001000110010110;
12'b000101110110: dataB <= 32'b10101111110011110010111100101111;
12'b000101110111: dataB <= 32'b00001110001011101101000111110100;
12'b000101111000: dataB <= 32'b00011011111010010111101010101100;
12'b000101111001: dataB <= 32'b00001000000100011000011111001101;
12'b000101111010: dataB <= 32'b10101101000110001100111001101110;
12'b000101111011: dataB <= 32'b00001000111011100001010011000101;
12'b000101111100: dataB <= 32'b10010110010110111000100011110011;
12'b000101111101: dataB <= 32'b00001011111101101011010101001010;
12'b000101111110: dataB <= 32'b11001111001110111000110111001110;
12'b000101111111: dataB <= 32'b00001111001011100011100101101010;
12'b000110000000: dataB <= 32'b10010111011001001010100001010010;
12'b000110000001: dataB <= 32'b00001011110100100101011101111100;
12'b000110000010: dataB <= 32'b00101110111111101010011011001100;
12'b000110000011: dataB <= 32'b00001011001011011011001111100100;
12'b000110000100: dataB <= 32'b01101010111001111110111101001010;
12'b000110000101: dataB <= 32'b00000111100011000110101001111110;
12'b000110000110: dataB <= 32'b10010010001110100000010111000110;
12'b000110000111: dataB <= 32'b00001100001010010101100001010011;
12'b000110001000: dataB <= 32'b11100111000101100101000011011000;
12'b000110001001: dataB <= 32'b00000101010001001011001111000100;
12'b000110001010: dataB <= 32'b00101101001100101011100101100001;
12'b000110001011: dataB <= 32'b00001100101111100001101011001100;
12'b000110001100: dataB <= 32'b11101001101011000010101010001110;
12'b000110001101: dataB <= 32'b00000111100110010001000011101101;
12'b000110001110: dataB <= 32'b01001110100100100100100000110000;
12'b000110001111: dataB <= 32'b00001110110000100011010100101011;
12'b000110010000: dataB <= 32'b00100110011101111000010011101011;
12'b000110010001: dataB <= 32'b00001001110000011111001100110110;
12'b000110010010: dataB <= 32'b11100101011010010001100010010100;
12'b000110010011: dataB <= 32'b00000111101000011010000111011010;
12'b000110010100: dataB <= 32'b10010110101001100011110011110011;
12'b000110010101: dataB <= 32'b00000000110100000011001001111001;
12'b000110010110: dataB <= 32'b01100110110010000000110101000010;
12'b000110010111: dataB <= 32'b00000111111110100001000001011111;
12'b000110011000: dataB <= 32'b01010001011101100010100011101100;
12'b000110011001: dataB <= 32'b00000001110010001100011011010001;
12'b000110011010: dataB <= 32'b00000110111100111100100000110001;
12'b000110011011: dataB <= 32'b00001100110001011111011100001101;
12'b000110011100: dataB <= 32'b11011100001110011100110101011100;
12'b000110011101: dataB <= 32'b00000110011000100010110101110010;
12'b000110011110: dataB <= 32'b00000101010111110011100110111110;
12'b000110011111: dataB <= 32'b00001011001100100100111101000100;
12'b000110100000: dataB <= 32'b11001101100110011001110011110101;
12'b000110100001: dataB <= 32'b00001000001011010011001110010010;
12'b000110100010: dataB <= 32'b01100011001010000111100111011010;
12'b000110100011: dataB <= 32'b00001110110110101111011111101010;
12'b000110100100: dataB <= 32'b00010100001001010010100010001110;
12'b000110100101: dataB <= 32'b00000000110010011110000101000010;
12'b000110100110: dataB <= 32'b00000100110001001011100111000100;
12'b000110100111: dataB <= 32'b00001110001101011101101001000011;
12'b000110101000: dataB <= 32'b10100101000110101111011011011001;
12'b000110101001: dataB <= 32'b00001011001000100010110010101011;
12'b000110101010: dataB <= 32'b10100101011110011110101101101110;
12'b000110101011: dataB <= 32'b00000110100010010100011001101111;
12'b000110101100: dataB <= 32'b00000000000001001110000101110100;
12'b000110101101: dataB <= 32'b00000000000000000000000000000000;
12'b000110101110: dataB <= 32'b11010111110010101111100111111110;
12'b000110101111: dataB <= 32'b00001001101011011011011011000000;
12'b000110110000: dataB <= 32'b00000011000011101011011101010001;
12'b000110110001: dataB <= 32'b00000111100001010010010000100101;
12'b000110110010: dataB <= 32'b11110011101101100010000100001011;
12'b000110110011: dataB <= 32'b00001010100001100000100111100101;
12'b000110110100: dataB <= 32'b10011111011110111101111001010101;
12'b000110110101: dataB <= 32'b00000100101110001011001011011001;
12'b000110110110: dataB <= 32'b11000101011110000010000110101100;
12'b000110110111: dataB <= 32'b00001000111001011011111001111000;
12'b000110111000: dataB <= 32'b10100011000111010001011011001011;
12'b000110111001: dataB <= 32'b00001000101000001011101010101011;
12'b000110111010: dataB <= 32'b00011001000001001010100001101011;
12'b000110111011: dataB <= 32'b00000100010110011100010101111011;
12'b000110111100: dataB <= 32'b10111000111000110010100000101111;
12'b000110111101: dataB <= 32'b00001000100001010010111111101101;
12'b000110111110: dataB <= 32'b10101110110011001011001010001110;
12'b000110111111: dataB <= 32'b00000100111101100100100110101110;
12'b000111000000: dataB <= 32'b11001010011101011000010000110000;
12'b000111000001: dataB <= 32'b00000111100111100000000101010000;
12'b000111000010: dataB <= 32'b10011011101001100010000010100101;
12'b000111000011: dataB <= 32'b00000111001001001101001010000111;
12'b000111000100: dataB <= 32'b00100101010101111100001000101010;
12'b000111000101: dataB <= 32'b00001001100001001101100110101100;
12'b000111000110: dataB <= 32'b00000111100011110010111110000111;
12'b000111000111: dataB <= 32'b00000111101011100000011001101010;
12'b000111001000: dataB <= 32'b00100101101001011101001000001000;
12'b000111001001: dataB <= 32'b00000001010110000011000011000111;
12'b000111001010: dataB <= 32'b01101101001010101010000100011010;
12'b000111001011: dataB <= 32'b00001100100100100001000110100110;
12'b000111001100: dataB <= 32'b11110101101011101010001100101101;
12'b000111001101: dataB <= 32'b00001101101001101101000011110011;
12'b000111001110: dataB <= 32'b10100001111010101111101010001011;
12'b000111001111: dataB <= 32'b00000111000100010100100011010100;
12'b000111010000: dataB <= 32'b01101101000010001100111001101110;
12'b000111010001: dataB <= 32'b00001001111010100011010011001101;
12'b000111010010: dataB <= 32'b11010010011010100000010011110100;
12'b000111010011: dataB <= 32'b00001100111011101101010001000010;
12'b000111010100: dataB <= 32'b11001111010010101000010111001111;
12'b000111010101: dataB <= 32'b00001110101000100111100001100010;
12'b000111010110: dataB <= 32'b10011011011101000010110001010101;
12'b000111010111: dataB <= 32'b00001100010011101001011001111100;
12'b000111011000: dataB <= 32'b01101100110111100001111010101011;
12'b000111011001: dataB <= 32'b00001010101001011101001111100011;
12'b000111011010: dataB <= 32'b01101010110110001110111100101000;
12'b000111011011: dataB <= 32'b00000110100100000100110110001110;
12'b000111011100: dataB <= 32'b11001110010010001000010110000111;
12'b000111011101: dataB <= 32'b00001011101000011001100101010011;
12'b000111011110: dataB <= 32'b01100111000101101101010100011010;
12'b000111011111: dataB <= 32'b00000101010010001011010111001100;
12'b000111100000: dataB <= 32'b10101101001000101100000100100010;
12'b000111100001: dataB <= 32'b00001100101110100101101011001011;
12'b000111100010: dataB <= 32'b00101101100110110010011001101101;
12'b000111100011: dataB <= 32'b00000111000110010001000111110101;
12'b000111100100: dataB <= 32'b11001100101000101101000000110011;
12'b000111100101: dataB <= 32'b00001110101110100101010100100011;
12'b000111100110: dataB <= 32'b10100010011001100000010011001101;
12'b000111100111: dataB <= 32'b00001001101111100001001101000110;
12'b000111101000: dataB <= 32'b01100111010110000001100010110110;
12'b000111101001: dataB <= 32'b00000110101001010100001011010010;
12'b000111101010: dataB <= 32'b10010100101101100100000100010101;
12'b000111101011: dataB <= 32'b00000001110111000011010101110001;
12'b000111101100: dataB <= 32'b01100110110001101000110011100011;
12'b000111101101: dataB <= 32'b00001001011110100001000001110111;
12'b000111101110: dataB <= 32'b11010101100001011010110011001110;
12'b000111101111: dataB <= 32'b00000010010101001010100010111000;
12'b000111110000: dataB <= 32'b11000111001001000100110001010100;
12'b000111110001: dataB <= 32'b00001100101111100001011100011101;
12'b000111110010: dataB <= 32'b11011000001110011100110110111101;
12'b000111110011: dataB <= 32'b00000111011001100010110101101010;
12'b000111110100: dataB <= 32'b01000111100011110010111000011110;
12'b000111110101: dataB <= 32'b00001010101011100100111101000100;
12'b000111110110: dataB <= 32'b11010001101010001001100100110110;
12'b000111110111: dataB <= 32'b00000111101011010101010010001010;
12'b000111111000: dataB <= 32'b11100101001010011111101000111010;
12'b000111111001: dataB <= 32'b00001111010011110011011011100001;
12'b000111111010: dataB <= 32'b01001110001101001010110010010000;
12'b000111111011: dataB <= 32'b00000001010101011000000100110010;
12'b000111111100: dataB <= 32'b01000010111101001011110101100100;
12'b000111111101: dataB <= 32'b00001101101010100001101001000011;
12'b000111111110: dataB <= 32'b01100101000111000111001100010111;
12'b000111111111: dataB <= 32'b00001010000111100010110010101011;
12'b001000000000: dataB <= 32'b10101001011010101110011101101011;
12'b001000000001: dataB <= 32'b00000101100011010010011101111111;
12'b001000000010: dataB <= 32'b00000000000001010110010110010100;
12'b001000000011: dataB <= 32'b00000000000000000000000000000000;
12'b001000000100: dataB <= 32'b10011101110110111111001001011110;
12'b001000000101: dataB <= 32'b00001001001010011101011010110000;
12'b001000000110: dataB <= 32'b10000011001111101010101101001111;
12'b001000000111: dataB <= 32'b00000110000001001110011000101101;
12'b001000001000: dataB <= 32'b01110111100101010010010011101101;
12'b001000001001: dataB <= 32'b00001001000001011100100111110101;
12'b001000001010: dataB <= 32'b00100001011111000101011001110100;
12'b001000001011: dataB <= 32'b00000100110000001101010011001001;
12'b001000001100: dataB <= 32'b11001001100101111010000110001100;
12'b001000001101: dataB <= 32'b00001001111000100001111001101000;
12'b001000001110: dataB <= 32'b01100011000110111000111010101010;
12'b001000001111: dataB <= 32'b00001000001000010001110010100011;
12'b001000010000: dataB <= 32'b00011001000101000010110001001110;
12'b001000010001: dataB <= 32'b00000100110111011000010101110011;
12'b001000010010: dataB <= 32'b11110110110000101011000000110001;
12'b001000010011: dataB <= 32'b00000111000001010011000111110100;
12'b001000010100: dataB <= 32'b01101100101011001010101001101110;
12'b001000010101: dataB <= 32'b00000110011110100010100110111110;
12'b001000010110: dataB <= 32'b01001000100101000000100000110010;
12'b001000010111: dataB <= 32'b00000111001000011010000100111001;
12'b001000011000: dataB <= 32'b10011111101001010010010001100111;
12'b001000011001: dataB <= 32'b00000110101010001111010010011111;
12'b001000011010: dataB <= 32'b11100111010001111100001000001001;
12'b001000011011: dataB <= 32'b00001000000001010001101110101011;
12'b001000011100: dataB <= 32'b01001011101011101010001101000100;
12'b001000011101: dataB <= 32'b00000111001011011100011001011010;
12'b001000011110: dataB <= 32'b10101001100101100101010111101000;
12'b001000011111: dataB <= 32'b00000010011001000011001011011110;
12'b001000100000: dataB <= 32'b00101101000110011001110101111100;
12'b001000100001: dataB <= 32'b00001011100010100001000110101110;
12'b001000100010: dataB <= 32'b00111001100011011001101100001011;
12'b001000100011: dataB <= 32'b00001100100111101100111011110011;
12'b001000100100: dataB <= 32'b00100111111010111111001001101010;
12'b001000100101: dataB <= 32'b00000101100101010010100111010100;
12'b001000100110: dataB <= 32'b11101100111010010100101001001101;
12'b001000100111: dataB <= 32'b00001010111001100011001111010100;
12'b001000101000: dataB <= 32'b01001110100010001000010100010110;
12'b001000101001: dataB <= 32'b00001101111001101111001100111011;
12'b001000101010: dataB <= 32'b00010001011010010000010111001111;
12'b001000101011: dataB <= 32'b00001101100110101001011101011011;
12'b001000101100: dataB <= 32'b10011101011100111011010010010111;
12'b001000101101: dataB <= 32'b00001100010001101011010110000100;
12'b001000101110: dataB <= 32'b11101100110011010001001010001010;
12'b001000101111: dataB <= 32'b00001010001000011101001111011010;
12'b001000110000: dataB <= 32'b01101000110010100110101011100110;
12'b001000110001: dataB <= 32'b00000101000101000101000010011110;
12'b001000110010: dataB <= 32'b00001010011001110000010101101000;
12'b001000110011: dataB <= 32'b00001010100111011101100101010100;
12'b001000110100: dataB <= 32'b11101001000001110101010101011011;
12'b001000110101: dataB <= 32'b00000101110011001111011111001011;
12'b001000110110: dataB <= 32'b00101101000100101100100011000100;
12'b001000110111: dataB <= 32'b00001100001100101001100111001011;
12'b001000111000: dataB <= 32'b01110001011110101010001001101100;
12'b001000111001: dataB <= 32'b00000110000111010001001111110100;
12'b001000111010: dataB <= 32'b01001010110000110101100001010110;
12'b001000111011: dataB <= 32'b00001110001011100111010000100100;
12'b001000111100: dataB <= 32'b11011110011001001000100010101111;
12'b001000111101: dataB <= 32'b00001001101110100011001101010110;
12'b001000111110: dataB <= 32'b11101001010001110001100011111000;
12'b001000111111: dataB <= 32'b00000110001001001110001111000001;
12'b001001000000: dataB <= 32'b11010010110101100100010100110110;
12'b001001000001: dataB <= 32'b00000010011001000111011101100001;
12'b001001000010: dataB <= 32'b01100100101101011001000010100101;
12'b001001000011: dataB <= 32'b00001010111110100001000010001111;
12'b001001000100: dataB <= 32'b01011001100101010011000011010000;
12'b001001000101: dataB <= 32'b00000010110111000110101110101000;
12'b001001000110: dataB <= 32'b01001001010001001101010001110110;
12'b001001000111: dataB <= 32'b00001100101101100101011000100110;
12'b001001001000: dataB <= 32'b11010100010010100100101000011101;
12'b001001001001: dataB <= 32'b00001000011001100000110101101010;
12'b001001001010: dataB <= 32'b11001011101011101010001001111110;
12'b001001001011: dataB <= 32'b00001010001010100100111001000100;
12'b001001001100: dataB <= 32'b10010111110001111001100101010111;
12'b001001001101: dataB <= 32'b00000111001011010111010110000010;
12'b001001001110: dataB <= 32'b00100101000110101111011001111010;
12'b001001001111: dataB <= 32'b00001111010000110101010011010001;
12'b001001010000: dataB <= 32'b11001010010101000011000010010010;
12'b001001010001: dataB <= 32'b00000001111000010010001000101010;
12'b001001010010: dataB <= 32'b11000011000101001100010100100101;
12'b001001010011: dataB <= 32'b00001101001000100101101000111011;
12'b001001010100: dataB <= 32'b00100101000011010110101100110110;
12'b001001010101: dataB <= 32'b00001001000110100000101110100011;
12'b001001010110: dataB <= 32'b10101011010110110110001101001001;
12'b001001010111: dataB <= 32'b00000100100100001110100110010111;
12'b001001011000: dataB <= 32'b00000000000001100110100110110101;
12'b001001011001: dataB <= 32'b00000000000000000000000000000000;
12'b001001011010: dataB <= 32'b01100001110111010110101010011110;
12'b001001011011: dataB <= 32'b00001000101010100001011110011000;
12'b001001011100: dataB <= 32'b00000101011011011010001101001100;
12'b001001011101: dataB <= 32'b00000100100010001010011100111110;
12'b001001011110: dataB <= 32'b10111011011001001010100011101111;
12'b001001011111: dataB <= 32'b00000111100001011010100111110100;
12'b001001100000: dataB <= 32'b10100101011111001100111010010011;
12'b001001100001: dataB <= 32'b00000100110001001111011010110000;
12'b001001100010: dataB <= 32'b00001101101101101010000110001101;
12'b001001100011: dataB <= 32'b00001010110111100111111001011001;
12'b001001100100: dataB <= 32'b00100011000110101000011010001001;
12'b001001100101: dataB <= 32'b00000111001000010101111010100011;
12'b001001100110: dataB <= 32'b00011001000101000011010001010000;
12'b001001100111: dataB <= 32'b00000101111000010100011001110011;
12'b001001101000: dataB <= 32'b00110100101000101011100001010100;
12'b001001101001: dataB <= 32'b00000101100001010011001011110100;
12'b001001101010: dataB <= 32'b11101010100110111010001001101101;
12'b001001101011: dataB <= 32'b00000111111110011110100011001101;
12'b001001101100: dataB <= 32'b10000110101100110001000001010101;
12'b001001101101: dataB <= 32'b00000110001000010110000100101001;
12'b001001101110: dataB <= 32'b01100101101001001010100001001001;
12'b001001101111: dataB <= 32'b00000110001010010001011010110111;
12'b001001110000: dataB <= 32'b10101001001101111100000111101001;
12'b001001110001: dataB <= 32'b00000110100001010101110010101011;
12'b001001110010: dataB <= 32'b10001111110011011001101011100011;
12'b001001110011: dataB <= 32'b00000110101011011000011001010010;
12'b001001110100: dataB <= 32'b11101101100001101101010110101000;
12'b001001110101: dataB <= 32'b00000010111011000101010111100101;
12'b001001110110: dataB <= 32'b10101110111110001001110110111100;
12'b001001110111: dataB <= 32'b00001010000001100001000110111101;
12'b001001111000: dataB <= 32'b01111011011011001001001011101001;
12'b001001111001: dataB <= 32'b00001100000101101100110111101010;
12'b001001111010: dataB <= 32'b01101101110111010110101001001010;
12'b001001111011: dataB <= 32'b00000100100110010000101111010011;
12'b001001111100: dataB <= 32'b01101100110110010100101001001101;
12'b001001111101: dataB <= 32'b00001011111000100101001111010100;
12'b001001111110: dataB <= 32'b11001100101001110000010101010111;
12'b001001111111: dataB <= 32'b00001110110110101111000100111011;
12'b001010000000: dataB <= 32'b01010101011101111000010111001111;
12'b001010000001: dataB <= 32'b00001100100100101101011001011011;
12'b001010000010: dataB <= 32'b10100001100000111011110010111010;
12'b001010000011: dataB <= 32'b00001100101111101101010010000100;
12'b001010000100: dataB <= 32'b01101010101110111000111001101001;
12'b001010000101: dataB <= 32'b00001001001000011111001111010010;
12'b001010000110: dataB <= 32'b00100110101110110110011011000101;
12'b001010000111: dataB <= 32'b00000100000110000101001010101110;
12'b001010001000: dataB <= 32'b01000110100001011000010100101001;
12'b001010001001: dataB <= 32'b00001001100110100001101001010100;
12'b001010001010: dataB <= 32'b01101000111101111101010110011100;
12'b001010001011: dataB <= 32'b00000110010100010011100111001011;
12'b001010001100: dataB <= 32'b10101110111100110101000010000110;
12'b001010001101: dataB <= 32'b00001011101010101101100011000010;
12'b001010001110: dataB <= 32'b10110011010110011001111001001100;
12'b001010001111: dataB <= 32'b00000101001000010011010011110011;
12'b001010010000: dataB <= 32'b11001010111001000110000001111000;
12'b001010010001: dataB <= 32'b00001101101001101001001100101100;
12'b001010010010: dataB <= 32'b00011010011000111001000010110001;
12'b001010010011: dataB <= 32'b00001001101110100011001101100111;
12'b001010010100: dataB <= 32'b01101011001101100001100100011010;
12'b001010010101: dataB <= 32'b00000101101010001010010110111001;
12'b001010010110: dataB <= 32'b00010010111001100100010101110111;
12'b001010010111: dataB <= 32'b00000011011011001011101001010010;
12'b001010011000: dataB <= 32'b01100010101101001001010001100111;
12'b001010011001: dataB <= 32'b00001011111100100001000010011111;
12'b001010011010: dataB <= 32'b01011101100101010011010011010010;
12'b001010011011: dataB <= 32'b00000011111001000110110110010000;
12'b001010011100: dataB <= 32'b11001011011001010101100010111000;
12'b001010011101: dataB <= 32'b00001100001011100111011000110110;
12'b001010011110: dataB <= 32'b00001110011010100100011001011101;
12'b001010011111: dataB <= 32'b00001001011001100000110101100011;
12'b001010100000: dataB <= 32'b00001111110011011001101011011101;
12'b001010100001: dataB <= 32'b00001001101001100100111001001101;
12'b001010100010: dataB <= 32'b10011011110001101001100110011000;
12'b001010100011: dataB <= 32'b00000110101011011001011001111010;
12'b001010100100: dataB <= 32'b11100101000111000111001010111001;
12'b001010100101: dataB <= 32'b00001111001101110101001010111000;
12'b001010100110: dataB <= 32'b01000110011101000011100010110100;
12'b001010100111: dataB <= 32'b00000010111010001110001100101011;
12'b001010101000: dataB <= 32'b01000101010001001100100011100111;
12'b001010101001: dataB <= 32'b00001100000110101001100100111100;
12'b001010101010: dataB <= 32'b11100101000011100110001101010100;
12'b001010101011: dataB <= 32'b00001000000110011110101110011010;
12'b001010101100: dataB <= 32'b01101101010011000101101100000111;
12'b001010101101: dataB <= 32'b00000011000110001100101110101111;
12'b001010101110: dataB <= 32'b00000000000001110110100111010101;
12'b001010101111: dataB <= 32'b00000000000000000000000000000000;
12'b001010110000: dataB <= 32'b00111010111111010001011111001011;
12'b001010110001: dataB <= 32'b00000101001110101110111100001011;
12'b001010110010: dataB <= 32'b00101101110101000001000110000101;
12'b001010110011: dataB <= 32'b00000001010110001111101011000110;
12'b001010110100: dataB <= 32'b01101100001001010101100111111000;
12'b001010110101: dataB <= 32'b00000000110000010011001010010000;
12'b001010110110: dataB <= 32'b01101110110110011001101001101011;
12'b001010110111: dataB <= 32'b00001000110110101101100000010010;
12'b001010111000: dataB <= 32'b00110111100101000100100110110011;
12'b001010111001: dataB <= 32'b00001011101010111100110000100101;
12'b001010111010: dataB <= 32'b11100010111000001010100100101011;
12'b001010111011: dataB <= 32'b00000100010001111101010101100010;
12'b001010111100: dataB <= 32'b01100011001101101101111000011101;
12'b001010111101: dataB <= 32'b00001100010100001101010101100100;
12'b001010111110: dataB <= 32'b01010100010101110110101010011101;
12'b001010111111: dataB <= 32'b00000000110100100101011010000000;
12'b001011000000: dataB <= 32'b10010010101001000010000110101100;
12'b001011000001: dataB <= 32'b00001111010000010001000010111001;
12'b001011000010: dataB <= 32'b10010111110000100110011010111101;
12'b001011000011: dataB <= 32'b00000100010011000011010000110110;
12'b001011000100: dataB <= 32'b01110100110101010101100100111101;
12'b001011000101: dataB <= 32'b00000101010011101101011111101010;
12'b001011000110: dataB <= 32'b10100110101110000100000100110000;
12'b001011000111: dataB <= 32'b00000000110010111001010101110010;
12'b001011001000: dataB <= 32'b01111001100000110001000001101000;
12'b001011001001: dataB <= 32'b00000101110010001101001101010101;
12'b001011001010: dataB <= 32'b11110000100110101100100100010010;
12'b001011001011: dataB <= 32'b00001101111010101011110110111000;
12'b001011001100: dataB <= 32'b00011110100000111011101110010010;
12'b001011001101: dataB <= 32'b00000000101011100010111110110010;
12'b001011001110: dataB <= 32'b10101100001000100001100100101000;
12'b001011001111: dataB <= 32'b00000010100111011010100101001000;
12'b001011010000: dataB <= 32'b01111010100111010001010101001101;
12'b001011010001: dataB <= 32'b00000011010110010111011101101001;
12'b001011010010: dataB <= 32'b01011010100110010011010110101101;
12'b001011010011: dataB <= 32'b00001100001000100110110110001001;
12'b001011010100: dataB <= 32'b00010101100100001100011011110101;
12'b001011010101: dataB <= 32'b00001011000010100010100001111110;
12'b001011010110: dataB <= 32'b00101111010100001100000111110001;
12'b001011010111: dataB <= 32'b00000010000110101100100101101101;
12'b001011011000: dataB <= 32'b11110000111101111110001101011010;
12'b001011011001: dataB <= 32'b00000111100110101000100110010011;
12'b001011011010: dataB <= 32'b01010110101000011010000100101100;
12'b001011011011: dataB <= 32'b00000100001101100111000001001001;
12'b001011011100: dataB <= 32'b10010110110011001010010010101001;
12'b001011011101: dataB <= 32'b00000011010111100101110111000010;
12'b001011011110: dataB <= 32'b01010001110000001101000100110110;
12'b001011011111: dataB <= 32'b00000011001100110100111110001101;
12'b001011100000: dataB <= 32'b10011110101110101100001110010011;
12'b001011100001: dataB <= 32'b00001010010011110011011001101001;
12'b001011100010: dataB <= 32'b11011110100010100110010011011011;
12'b001011100011: dataB <= 32'b00000101001000110000100101010001;
12'b001011100100: dataB <= 32'b01101010011000111011000110001101;
12'b001011100101: dataB <= 32'b00000100010101101001011001110000;
12'b001011100110: dataB <= 32'b10011101101011000101111100011100;
12'b001011100111: dataB <= 32'b00000100100100100110101110011110;
12'b001011101000: dataB <= 32'b11001101001000100110001000111010;
12'b001011101001: dataB <= 32'b00000111001100100110111011100100;
12'b001011101010: dataB <= 32'b00100110101000110100111101010111;
12'b001011101011: dataB <= 32'b00000101010100001011101000101010;
12'b001011101100: dataB <= 32'b01011101011010001100111011110100;
12'b001011101101: dataB <= 32'b00001101111001110101101001000101;
12'b001011101110: dataB <= 32'b00010110111000101101100011111100;
12'b001011101111: dataB <= 32'b00001110001000100000111111101011;
12'b001011110000: dataB <= 32'b01110011000101101101011001011001;
12'b001011110001: dataB <= 32'b00001100111000011011110000001011;
12'b001011110010: dataB <= 32'b01101101101010110101011100011010;
12'b001011110011: dataB <= 32'b00000101100111101100110011011110;
12'b001011110100: dataB <= 32'b11001101100010001010111110101101;
12'b001011110101: dataB <= 32'b00001100101101011010111101100100;
12'b001011110110: dataB <= 32'b10111001100000110001001110101001;
12'b001011110111: dataB <= 32'b00000100101100011100110110100101;
12'b001011111000: dataB <= 32'b00111001001000110100101100010011;
12'b001011111001: dataB <= 32'b00000101110010101101001101010100;
12'b001011111010: dataB <= 32'b00100010110111100001111100101010;
12'b001011111011: dataB <= 32'b00000110100001100100010100011010;
12'b001011111100: dataB <= 32'b10001111110001110101111010011010;
12'b001011111101: dataB <= 32'b00001101011010000111100001101110;
12'b001011111110: dataB <= 32'b00101001110110010101100011111000;
12'b001011111111: dataB <= 32'b00000011000111110010101110001110;
12'b001100000000: dataB <= 32'b00100000110111000000111010000101;
12'b001100000001: dataB <= 32'b00000011001111010111000001011011;
12'b001100000010: dataB <= 32'b10101000100110110001110011100111;
12'b001100000011: dataB <= 32'b00000011011001010111100111101010;
12'b001100000100: dataB <= 32'b00000000000011010100011010110001;
12'b001100000101: dataB <= 32'b00000000000000000000000000000000;
12'b001100000110: dataB <= 32'b01111011000111100010001111001101;
12'b001100000111: dataB <= 32'b00000101001101101101000100010010;
12'b001100001000: dataB <= 32'b10100111111001010000100111100101;
12'b001100001001: dataB <= 32'b00000000110011001101100010110110;
12'b001100001010: dataB <= 32'b01110010010001001101010110111000;
12'b001100001011: dataB <= 32'b00000000101101010011000110101000;
12'b001100001100: dataB <= 32'b10101110111110101001111010001100;
12'b001100001101: dataB <= 32'b00001000010110101001100100100001;
12'b001100001110: dataB <= 32'b10110011101101000100000110010011;
12'b001100001111: dataB <= 32'b00001100001100111100111100011100;
12'b001100010000: dataB <= 32'b11100010111000011010000101001010;
12'b001100010001: dataB <= 32'b00000100001111111001011101101010;
12'b001100010010: dataB <= 32'b01100011001101011101110111011101;
12'b001100010011: dataB <= 32'b00001011110110001011001101100100;
12'b001100010100: dataB <= 32'b01011000010001100110101000111110;
12'b001100010101: dataB <= 32'b00000000110001100011011010011000;
12'b001100010110: dataB <= 32'b00010100100101010001100111001100;
12'b001100010111: dataB <= 32'b00001111010011010010111011001010;
12'b001100011000: dataB <= 32'b00010011101100010101111001011110;
12'b001100011001: dataB <= 32'b00000100010001000011001000101110;
12'b001100011010: dataB <= 32'b00110101000001001101010011111100;
12'b001100011011: dataB <= 32'b00000101010010101001100011110011;
12'b001100011100: dataB <= 32'b10101000110010000100000100101111;
12'b001100011101: dataB <= 32'b00000000101111110111011101111010;
12'b001100011110: dataB <= 32'b00110101101001000000100010000101;
12'b001100011111: dataB <= 32'b00000101110001001101000101001101;
12'b001100100000: dataB <= 32'b00110010101110101100110100010000;
12'b001100100001: dataB <= 32'b00001100111011100101111011010001;
12'b001100100010: dataB <= 32'b10100010100100111011001110010100;
12'b001100100011: dataB <= 32'b00000001001000100010111111000010;
12'b001100100100: dataB <= 32'b01110000001100110001000101100111;
12'b001100100101: dataB <= 32'b00000011100110011100100101100000;
12'b001100100110: dataB <= 32'b01111100110011100010000101001100;
12'b001100100111: dataB <= 32'b00000010110100010011011010000001;
12'b001100101000: dataB <= 32'b01011100100110010011010110101101;
12'b001100101001: dataB <= 32'b00001100101010100110111010011001;
12'b001100101010: dataB <= 32'b00010001100000001011101011010111;
12'b001100101011: dataB <= 32'b00001100100100100110100001101110;
12'b001100101100: dataB <= 32'b00101101011100001011010111110001;
12'b001100101101: dataB <= 32'b00000011000100101110101101100101;
12'b001100101110: dataB <= 32'b11101111000101101110001011111011;
12'b001100101111: dataB <= 32'b00001000100111101010101010010011;
12'b001100110000: dataB <= 32'b00011000100100100001010101001011;
12'b001100110001: dataB <= 32'b00000100001011100111000101011001;
12'b001100110010: dataB <= 32'b00011000101111010010110011001000;
12'b001100110011: dataB <= 32'b00000010110101100001110111001011;
12'b001100110100: dataB <= 32'b01001101101000001100010100010100;
12'b001100110101: dataB <= 32'b00000011101010110011000110000101;
12'b001100110110: dataB <= 32'b10100000101110101100011101110101;
12'b001100110111: dataB <= 32'b00001001110100101111100001111001;
12'b001100111000: dataB <= 32'b10100010100110010110100010011001;
12'b001100111001: dataB <= 32'b00000110000111110010101101100001;
12'b001100111010: dataB <= 32'b01101110011101000010100110001100;
12'b001100111011: dataB <= 32'b00000011110011100111011110001000;
12'b001100111100: dataB <= 32'b11011001101010110110011011011101;
12'b001100111101: dataB <= 32'b00000101100011101000110010001110;
12'b001100111110: dataB <= 32'b01001101000000010101100111111010;
12'b001100111111: dataB <= 32'b00000111001100100110111011011101;
12'b001101000000: dataB <= 32'b11101000101100110100011100011000;
12'b001101000001: dataB <= 32'b00000100110011000111100000111001;
12'b001101000010: dataB <= 32'b11011011011010001100111011010110;
12'b001101000011: dataB <= 32'b00001100111011101111110000111100;
12'b001101000100: dataB <= 32'b10010110110100100101000010111010;
12'b001101000101: dataB <= 32'b00001111001010100000111111101011;
12'b001101000110: dataB <= 32'b10110011001101100101011000011001;
12'b001101000111: dataB <= 32'b00001011111010010111110000001010;
12'b001101001000: dataB <= 32'b11101001101110101101101011011100;
12'b001101001001: dataB <= 32'b00000110100110101100110111001110;
12'b001101001010: dataB <= 32'b10001001010110010010111110101111;
12'b001101001011: dataB <= 32'b00001100101111011010111101011100;
12'b001101001100: dataB <= 32'b11110101101001000000101111001100;
12'b001101001101: dataB <= 32'b00000101001011011100110110011101;
12'b001101001110: dataB <= 32'b11111001010000110100001011110101;
12'b001101001111: dataB <= 32'b00000101110001101011010001010011;
12'b001101010000: dataB <= 32'b01100010110111101010101101001100;
12'b001101010001: dataB <= 32'b00001000000001101000010100100001;
12'b001101010010: dataB <= 32'b10001011101001100101111001011011;
12'b001101010011: dataB <= 32'b00001100011100000101011001011110;
12'b001101010100: dataB <= 32'b00100011111010001101100010110110;
12'b001101010101: dataB <= 32'b00000100000101110100110101111110;
12'b001101010110: dataB <= 32'b11100000110111010001011011000110;
12'b001101010111: dataB <= 32'b00000011001101010110111101100010;
12'b001101011000: dataB <= 32'b01101010101011000010010100100101;
12'b001101011001: dataB <= 32'b00000010010110010011100011110011;
12'b001101011010: dataB <= 32'b00000000000011010100111010110010;
12'b001101011011: dataB <= 32'b00000000000000000000000000000000;
12'b001101011100: dataB <= 32'b11111001010011110010101111010000;
12'b001101011101: dataB <= 32'b00000101101100101101001000011001;
12'b001101011110: dataB <= 32'b11100001111001101000101000100101;
12'b001101011111: dataB <= 32'b00000000110000001001011010100110;
12'b001101100000: dataB <= 32'b11110110011001000100110101110111;
12'b001101100001: dataB <= 32'b00000000101010010010111110111000;
12'b001101100010: dataB <= 32'b00101111000010111010001010101101;
12'b001101100011: dataB <= 32'b00000111010110100101101000110001;
12'b001101100100: dataB <= 32'b00101111110101000011110110010010;
12'b001101100101: dataB <= 32'b00001100101110111101001000011100;
12'b001101100110: dataB <= 32'b10100010111000101001010101101001;
12'b001101100111: dataB <= 32'b00000100001110110101101001110010;
12'b001101101000: dataB <= 32'b00100001001101010101100101111100;
12'b001101101001: dataB <= 32'b00001011010111001011000101100100;
12'b001101101010: dataB <= 32'b10011100001101010110010111111110;
12'b001101101011: dataB <= 32'b00000000101110011111011010110000;
12'b001101101100: dataB <= 32'b10011000100001100001100111001011;
12'b001101101101: dataB <= 32'b00001110110110010010110111010010;
12'b001101101110: dataB <= 32'b01001111101000001101001000011110;
12'b001101101111: dataB <= 32'b00000011110000000010111100011101;
12'b001101110000: dataB <= 32'b11110101001001000100110010111010;
12'b001101110001: dataB <= 32'b00000100110001100101100111110011;
12'b001101110010: dataB <= 32'b10101010110110000100000101001110;
12'b001101110011: dataB <= 32'b00000000101100110011100110000010;
12'b001101110100: dataB <= 32'b10110001110001011000010011100011;
12'b001101110101: dataB <= 32'b00000101110000001100111101000100;
12'b001101110110: dataB <= 32'b11110100110110100101000100001111;
12'b001101110111: dataB <= 32'b00001011011101100001111011100001;
12'b001101111000: dataB <= 32'b11100100100101000010101101010111;
12'b001101111001: dataB <= 32'b00000010000110100010111111001010;
12'b001101111010: dataB <= 32'b01110100010101000000100110100110;
12'b001101111011: dataB <= 32'b00000100100100100000100101111000;
12'b001101111100: dataB <= 32'b01111100111111110010100101101011;
12'b001101111101: dataB <= 32'b00000010010001010001010110010001;
12'b001101111110: dataB <= 32'b10100000100110011011100111001100;
12'b001101111111: dataB <= 32'b00001101001100101000111010101001;
12'b001110000000: dataB <= 32'b11001101011000001010111010011000;
12'b001110000001: dataB <= 32'b00001101100110101000100101011101;
12'b001110000010: dataB <= 32'b11101001100000001010100111110001;
12'b001110000011: dataB <= 32'b00000100000010110000110001011100;
12'b001110000100: dataB <= 32'b00101111001001011101111010111101;
12'b001110000101: dataB <= 32'b00001001100111101100101110010100;
12'b001110000110: dataB <= 32'b11011010100100111000110101101010;
12'b001110000111: dataB <= 32'b00000100101010100111000101101000;
12'b001110001000: dataB <= 32'b10011010101011011011100100000110;
12'b001110001001: dataB <= 32'b00000010010010011011110111001011;
12'b001110001010: dataB <= 32'b01001001100000001011100011110011;
12'b001110001011: dataB <= 32'b00000100001000110011001101111101;
12'b001110001100: dataB <= 32'b10100010110010101100101101010111;
12'b001110001101: dataB <= 32'b00001001010101101011101010001001;
12'b001110001110: dataB <= 32'b10100100100110000110100001010110;
12'b001110001111: dataB <= 32'b00000111000110110100110101110001;
12'b001110010000: dataB <= 32'b01110010100101001010010110101100;
12'b001110010001: dataB <= 32'b00000011010001100011011110100000;
12'b001110010010: dataB <= 32'b11010101100110100110101001111110;
12'b001110010011: dataB <= 32'b00000111000010101010110101111110;
12'b001110010100: dataB <= 32'b11001100111000001100110110111001;
12'b001110010101: dataB <= 32'b00000111101100100110111111010101;
12'b001110010110: dataB <= 32'b01101010110000110011111011011010;
12'b001110010111: dataB <= 32'b00000100110010000101010101001001;
12'b001110011000: dataB <= 32'b01010111010110000100111010110111;
12'b001110011001: dataB <= 32'b00001011111100101011111000110100;
12'b001110011010: dataB <= 32'b01011000110000011100100001111000;
12'b001110011011: dataB <= 32'b00001111001101100000111111101100;
12'b001110011100: dataB <= 32'b00110001010101011101000111011001;
12'b001110011101: dataB <= 32'b00001010111011010001101000011010;
12'b001110011110: dataB <= 32'b00100101110010011101111010011101;
12'b001110011111: dataB <= 32'b00000111100110101110111110111111;
12'b001110100000: dataB <= 32'b10000111001110011011001110110010;
12'b001110100001: dataB <= 32'b00001100110001011010111001011100;
12'b001110100010: dataB <= 32'b11110001110001011000011111001111;
12'b001110100011: dataB <= 32'b00000101101010011110110110001101;
12'b001110100100: dataB <= 32'b10110101011100110011101011010110;
12'b001110100101: dataB <= 32'b00000101110000101001010101011011;
12'b001110100110: dataB <= 32'b11100100110111110011001101001110;
12'b001110100111: dataB <= 32'b00001001100001101100011000111000;
12'b001110101000: dataB <= 32'b01000111100001011101101000011011;
12'b001110101001: dataB <= 32'b00001010111101000011001101001110;
12'b001110101010: dataB <= 32'b11011111111001111101100010010100;
12'b001110101011: dataB <= 32'b00000101000100110100111101101101;
12'b001110101100: dataB <= 32'b10100010110111100001111011100111;
12'b001110101101: dataB <= 32'b00000011101011011000111001101010;
12'b001110101110: dataB <= 32'b00101100101111001010100101100100;
12'b001110101111: dataB <= 32'b00000001110100001111011011110100;
12'b001110110000: dataB <= 32'b00000000000011001101011010010011;
12'b001110110001: dataB <= 32'b00000000000000000000000000000000;
12'b001110110010: dataB <= 32'b01110111011011110011011111010011;
12'b001110110011: dataB <= 32'b00000101101011101101001100101001;
12'b001110110100: dataB <= 32'b11011011111010000000011001100101;
12'b001110110101: dataB <= 32'b00000000101101000111010010001110;
12'b001110110110: dataB <= 32'b01111010100000111100100101010110;
12'b001110110111: dataB <= 32'b00000001101000010010111011010001;
12'b001110111000: dataB <= 32'b10101111001011000010101010101110;
12'b001110111001: dataB <= 32'b00000110110101100001101001000000;
12'b001110111010: dataB <= 32'b01101001111001000011010101110001;
12'b001110111011: dataB <= 32'b00001100101111111101010100011011;
12'b001110111100: dataB <= 32'b10100100111100111000110110101000;
12'b001110111101: dataB <= 32'b00000100101101110001110001111010;
12'b001110111110: dataB <= 32'b11011111001101001101000100111011;
12'b001110111111: dataB <= 32'b00001010011000001010111001100011;
12'b001111000000: dataB <= 32'b11100000001101001110000110011101;
12'b001111000001: dataB <= 32'b00000000101011011101011011000000;
12'b001111000010: dataB <= 32'b00011010011101110001010111101011;
12'b001111000011: dataB <= 32'b00001110011000010010110011011011;
12'b001111000100: dataB <= 32'b11001011100000001100010110111110;
12'b001111000101: dataB <= 32'b00000100001110000010110000010100;
12'b001111000110: dataB <= 32'b10110011010000111100100001110111;
12'b001111000111: dataB <= 32'b00000100101111100001100111110100;
12'b001111001000: dataB <= 32'b10101010111010000100000101001100;
12'b001111001001: dataB <= 32'b00000001001001101111101110001010;
12'b001111001010: dataB <= 32'b01101011110101110000010100100010;
12'b001111001011: dataB <= 32'b00000101101111001100110101000100;
12'b001111001100: dataB <= 32'b01110100111110011101010100001101;
12'b001111001101: dataB <= 32'b00001001111110011011111011101010;
12'b001111001110: dataB <= 32'b01100110100101001010011100111001;
12'b001111001111: dataB <= 32'b00000011000100100010111111001011;
12'b001111010000: dataB <= 32'b01111000100001011000010111100110;
12'b001111010001: dataB <= 32'b00000101100011100010100110010000;
12'b001111010010: dataB <= 32'b10111101001011110011010110001010;
12'b001111010011: dataB <= 32'b00000010001111001111001110100001;
12'b001111010100: dataB <= 32'b11100010100110011011100111001100;
12'b001111010101: dataB <= 32'b00001101101110101000111110110001;
12'b001111010110: dataB <= 32'b10001011010000010010001001111000;
12'b001111010111: dataB <= 32'b00001110101000101010101001010101;
12'b001111011000: dataB <= 32'b10100111100000011010000111010001;
12'b001111011001: dataB <= 32'b00000101100001110010111001011100;
12'b001111011010: dataB <= 32'b00101101010001010101101001011101;
12'b001111011011: dataB <= 32'b00001010001000101110110110010100;
12'b001111011100: dataB <= 32'b11011110100001001000100110001001;
12'b001111011101: dataB <= 32'b00000101101001100111001010000000;
12'b001111011110: dataB <= 32'b00011100101011011100000101000101;
12'b001111011111: dataB <= 32'b00000001110000010101110011001100;
12'b001111100000: dataB <= 32'b01000111011000001010110011010001;
12'b001111100001: dataB <= 32'b00000101000111110001010101110101;
12'b001111100010: dataB <= 32'b11100010110010100100111100011001;
12'b001111100011: dataB <= 32'b00001000110101100111101010011001;
12'b001111100100: dataB <= 32'b10100110100101110110100000110100;
12'b001111100101: dataB <= 32'b00000111100110110100111110000001;
12'b001111100110: dataB <= 32'b10110100101101010001110111001011;
12'b001111100111: dataB <= 32'b00000011010000100001011110111000;
12'b001111101000: dataB <= 32'b10010011100010010110111000011110;
12'b001111101001: dataB <= 32'b00001000000010101010111001101110;
12'b001111101010: dataB <= 32'b01001110110000001100000101111000;
12'b001111101011: dataB <= 32'b00001000001100100111000011000110;
12'b001111101100: dataB <= 32'b00101100110100110011011010011011;
12'b001111101101: dataB <= 32'b00000100010000000011001001011001;
12'b001111101110: dataB <= 32'b00010101010001111100111001111000;
12'b001111101111: dataB <= 32'b00001010011110100101111000110100;
12'b001111110000: dataB <= 32'b00011000110000011011110001010101;
12'b001111110001: dataB <= 32'b00001111010000100000111111101101;
12'b001111110010: dataB <= 32'b01101111011101010100110110011000;
12'b001111110011: dataB <= 32'b00001001011100001101100100101001;
12'b001111110100: dataB <= 32'b10011111110010010110001000111110;
12'b001111110101: dataB <= 32'b00001000100110101111000010100111;
12'b001111110110: dataB <= 32'b01000111000110011011001110010101;
12'b001111110111: dataB <= 32'b00001100010011011010111001011100;
12'b001111111000: dataB <= 32'b11101011110101110000011111010010;
12'b001111111001: dataB <= 32'b00000110001001011110110110000101;
12'b001111111010: dataB <= 32'b01110011100100111011001010111000;
12'b001111111011: dataB <= 32'b00000101101111100111011001011011;
12'b001111111100: dataB <= 32'b10100100111011110011111101010001;
12'b001111111101: dataB <= 32'b00001011000010101110100001001000;
12'b001111111110: dataB <= 32'b11000101010101010101010111011011;
12'b001111111111: dataB <= 32'b00001001011110000011000001000101;
12'b010000000000: dataB <= 32'b11011001110101110101100010010001;
12'b010000000001: dataB <= 32'b00000110100011110101000101100101;
12'b010000000010: dataB <= 32'b10100010110111101010101100101001;
12'b010000000011: dataB <= 32'b00000100001001011000111001110010;
12'b010000000100: dataB <= 32'b10101110110111010011000111000100;
12'b010000000101: dataB <= 32'b00000001010010001101010111110100;
12'b010000000110: dataB <= 32'b00000000000011000101101010010100;
12'b010000000111: dataB <= 32'b00000000000000000000000000000000;
12'b010000001000: dataB <= 32'b11110011100011110100001110110110;
12'b010000001001: dataB <= 32'b00000110001010101011010001000000;
12'b010000001010: dataB <= 32'b00010111111010010000101010100110;
12'b010000001011: dataB <= 32'b00000000101010000111000101111111;
12'b010000001100: dataB <= 32'b11111100101100111100000100110101;
12'b010000001101: dataB <= 32'b00000010100101010010110111100001;
12'b010000001110: dataB <= 32'b01101101001111001010111010101111;
12'b010000001111: dataB <= 32'b00000110010101011101101001011000;
12'b010000010000: dataB <= 32'b11100011111001001011000101110000;
12'b010000010001: dataB <= 32'b00001100110001111001011100100010;
12'b010000010010: dataB <= 32'b10100100111101001000100111001000;
12'b010000010011: dataB <= 32'b00000101001011101101110110000010;
12'b010000010100: dataB <= 32'b10011101001101000100110011111001;
12'b010000010101: dataB <= 32'b00001001011001001010110001100011;
12'b010000010110: dataB <= 32'b01100110010000111101100100111100;
12'b010000010111: dataB <= 32'b00000001001000011011011011010001;
12'b010000011000: dataB <= 32'b11011110011110000001011000001011;
12'b010000011001: dataB <= 32'b00001101011010010100101111100011;
12'b010000011010: dataB <= 32'b00001001010100001011100101011101;
12'b010000011011: dataB <= 32'b00000100001101000100100100010100;
12'b010000011100: dataB <= 32'b00110001010100111100000000110101;
12'b010000011101: dataB <= 32'b00000100101110011111100111110101;
12'b010000011110: dataB <= 32'b11101010111110000100000101101011;
12'b010000011111: dataB <= 32'b00000001100111101011110010010010;
12'b010000100000: dataB <= 32'b11100101111010001000010110000001;
12'b010000100001: dataB <= 32'b00000101101110001110101101000011;
12'b010000100010: dataB <= 32'b00110101000110010101010100101100;
12'b010000100011: dataB <= 32'b00001000011110010101110111110011;
12'b010000100100: dataB <= 32'b11101000101001011010001011111010;
12'b010000100101: dataB <= 32'b00000100000010100011000011001011;
12'b010000100110: dataB <= 32'b01111100101001110000011000000110;
12'b010000100111: dataB <= 32'b00000111000011100100100110101000;
12'b010000101000: dataB <= 32'b11111101010111110100000110101010;
12'b010000101001: dataB <= 32'b00000010001101001111000110101001;
12'b010000101010: dataB <= 32'b01100100100110011011110111101100;
12'b010000101011: dataB <= 32'b00001101110001101001000011000010;
12'b010000101100: dataB <= 32'b01001011001000100001101000111001;
12'b010000101101: dataB <= 32'b00001111001011101100101101001101;
12'b010000101110: dataB <= 32'b01100011100100101001010111010001;
12'b010000101111: dataB <= 32'b00000111000001110011000001010100;
12'b010000110000: dataB <= 32'b00101011010101001101011000011110;
12'b010000110001: dataB <= 32'b00001011001001101110111010010100;
12'b010000110010: dataB <= 32'b11100000100001100000010110101000;
12'b010000110011: dataB <= 32'b00000110001000100101001110010000;
12'b010000110100: dataB <= 32'b10011110101011011100100110000100;
12'b010000110101: dataB <= 32'b00000010001110010001101111001100;
12'b010000110110: dataB <= 32'b00000101001100010010000011001111;
12'b010000110111: dataB <= 32'b00000101100110101111011101101101;
12'b010000111000: dataB <= 32'b11100100110010011101001011011011;
12'b010000111001: dataB <= 32'b00001000010101100011101110101001;
12'b010000111010: dataB <= 32'b10101000101001100110010000110001;
12'b010000111011: dataB <= 32'b00001000100110110101000110010001;
12'b010000111100: dataB <= 32'b00110100110101100001110111101011;
12'b010000111101: dataB <= 32'b00000011001110011101011111001001;
12'b010000111110: dataB <= 32'b10001111011010000110110110111110;
12'b010000111111: dataB <= 32'b00001001100010101010111101011110;
12'b010001000000: dataB <= 32'b11001110101000001011010100110111;
12'b010001000001: dataB <= 32'b00001000101100100111000110110110;
12'b010001000010: dataB <= 32'b11101100111000111010111001011100;
12'b010001000011: dataB <= 32'b00000100001111000010111101101000;
12'b010001000100: dataB <= 32'b10010011001101110100111000111000;
12'b010001000101: dataB <= 32'b00001001011110011111111000110011;
12'b010001000110: dataB <= 32'b10011010101100011011010000110010;
12'b010001000111: dataB <= 32'b00001111010011100000111111100101;
12'b010001001000: dataB <= 32'b11101011100001010100100101011000;
12'b010001001001: dataB <= 32'b00001000011100001011011100111000;
12'b010001001010: dataB <= 32'b10011011110010000110000111011110;
12'b010001001011: dataB <= 32'b00001001100111101101001010010111;
12'b010001001100: dataB <= 32'b00000110111010100011011101110111;
12'b010001001101: dataB <= 32'b00001100010101011100110101011100;
12'b010001001110: dataB <= 32'b11100101111010001000011111010100;
12'b010001001111: dataB <= 32'b00000110101000100000110101110101;
12'b010001010000: dataB <= 32'b00101111101000111010101001111000;
12'b010001010001: dataB <= 32'b00000101101110100101011101100011;
12'b010001010010: dataB <= 32'b01100100111011110100101101010011;
12'b010001010011: dataB <= 32'b00001100000011110010100101100000;
12'b010001010100: dataB <= 32'b10000011001001001101000110011010;
12'b010001010101: dataB <= 32'b00000111111110000010110100110101;
12'b010001010110: dataB <= 32'b10010011110001101101100001101111;
12'b010001010111: dataB <= 32'b00000111100011110011001101011101;
12'b010001011000: dataB <= 32'b10100100111011110011011101001011;
12'b010001011001: dataB <= 32'b00000100101000011000110101111010;
12'b010001011010: dataB <= 32'b01101110111011010011101000000011;
12'b010001011011: dataB <= 32'b00000001001111001011001111101101;
12'b010001011100: dataB <= 32'b00000000000010110110001001110101;
12'b010001011101: dataB <= 32'b00000000000000000000000000000000;
12'b010001011110: dataB <= 32'b01101111101011110100111110011000;
12'b010001011111: dataB <= 32'b00000111001010101001010101010000;
12'b010001100000: dataB <= 32'b11010001110010101000101011000111;
12'b010001100001: dataB <= 32'b00000001101000000100111101101110;
12'b010001100010: dataB <= 32'b01111100111000111011100100010100;
12'b010001100011: dataB <= 32'b00000011100011010100110011101010;
12'b010001100100: dataB <= 32'b01101011010011010011011010110000;
12'b010001100101: dataB <= 32'b00000101110100011001100101110000;
12'b010001100110: dataB <= 32'b01011101111001010010110101110000;
12'b010001100111: dataB <= 32'b00001100010011110101101000101010;
12'b010001101000: dataB <= 32'b10100100111101100000011000000111;
12'b010001101001: dataB <= 32'b00000101001010100111111010001010;
12'b010001101010: dataB <= 32'b10011101001101000100100010110111;
12'b010001101011: dataB <= 32'b00001000011001001100101001100011;
12'b010001101100: dataB <= 32'b00101010010100110101010011111011;
12'b010001101101: dataB <= 32'b00000010000110011001010111100010;
12'b010001101110: dataB <= 32'b01100010011110010001011000101011;
12'b010001101111: dataB <= 32'b00001011111100010110101011100100;
12'b010001110000: dataB <= 32'b10000111001100001010110011111100;
12'b010001110001: dataB <= 32'b00000100101011000110011100010011;
12'b010001110010: dataB <= 32'b11101111011100111011100000110010;
12'b010001110011: dataB <= 32'b00000101001101011011100111100101;
12'b010001110100: dataB <= 32'b11101011000010000100000110001011;
12'b010001110101: dataB <= 32'b00000010100101100101110110011010;
12'b010001110110: dataB <= 32'b10011111111010100000010111100001;
12'b010001110111: dataB <= 32'b00000101101101010000100101000011;
12'b010001111000: dataB <= 32'b11110011001110001101100101001011;
12'b010001111001: dataB <= 32'b00000110111110001111110011110011;
12'b010001111010: dataB <= 32'b01101010101101100001111010111011;
12'b010001111011: dataB <= 32'b00000101100001100011000011001100;
12'b010001111100: dataB <= 32'b11111100110110001000011001000110;
12'b010001111101: dataB <= 32'b00001000000010100110101010111000;
12'b010001111110: dataB <= 32'b00111001011111110100110111001001;
12'b010001111111: dataB <= 32'b00000010101011001111000010111010;
12'b010010000000: dataB <= 32'b10100110101010011100001000001100;
12'b010010000001: dataB <= 32'b00001101010011101001000111001010;
12'b010010000010: dataB <= 32'b00001001000000110001000111111001;
12'b010010000011: dataB <= 32'b00001111001110101110110101000101;
12'b010010000100: dataB <= 32'b00011111100100111000110111010000;
12'b010010000101: dataB <= 32'b00001000100001110011000101010100;
12'b010010000110: dataB <= 32'b01101001011001000101000110111101;
12'b010010000111: dataB <= 32'b00001011101010110001000010001100;
12'b010010001000: dataB <= 32'b00100100100101111000010111101000;
12'b010010001001: dataB <= 32'b00000110101000100011001110101001;
12'b010010001010: dataB <= 32'b00100000101011010101000111100011;
12'b010010001011: dataB <= 32'b00000010001011001101100111001101;
12'b010010001100: dataB <= 32'b00000011000000100001100011001110;
12'b010010001101: dataB <= 32'b00000110100101101011100001100101;
12'b010010001110: dataB <= 32'b01100110110110010101011010011100;
12'b010010001111: dataB <= 32'b00000111110101011111101110110010;
12'b010010010000: dataB <= 32'b10101010101101010110000000101110;
12'b010010010001: dataB <= 32'b00001001100111110011001110100001;
12'b010010010010: dataB <= 32'b10110110111101110001100111101011;
12'b010010010011: dataB <= 32'b00000011101100011011011111011001;
12'b010010010100: dataB <= 32'b01001101010101110110110101011110;
12'b010010010101: dataB <= 32'b00001010100011101011000001001110;
12'b010010010110: dataB <= 32'b00010010100100001010110100010110;
12'b010010010111: dataB <= 32'b00001000101100100111000110100111;
12'b010010011000: dataB <= 32'b11101100111101000010010111111100;
12'b010010011001: dataB <= 32'b00000100101101000010110010000000;
12'b010010011010: dataB <= 32'b00010011001001110100111000011000;
12'b010010011011: dataB <= 32'b00000111111110011001111000111011;
12'b010010011100: dataB <= 32'b01011100101100100010100000101111;
12'b010010011101: dataB <= 32'b00001110110110100000111111010110;
12'b010010011110: dataB <= 32'b10100111100101001100010100110110;
12'b010010011111: dataB <= 32'b00000110111100001001010101001000;
12'b010010100000: dataB <= 32'b10010101101101110110000101111101;
12'b010010100001: dataB <= 32'b00001010000111101101001101111111;
12'b010010100010: dataB <= 32'b11000110110010100011101100111001;
12'b010010100011: dataB <= 32'b00001011010110011100110101011011;
12'b010010100100: dataB <= 32'b11100001111010100000011110010111;
12'b010010100101: dataB <= 32'b00000111101000100000110101101101;
12'b010010100110: dataB <= 32'b00101011101101001010011000111001;
12'b010010100111: dataB <= 32'b00000101101101100001011101100011;
12'b010010101000: dataB <= 32'b01100110111111101101011100110101;
12'b010010101001: dataB <= 32'b00001101000101110100101101111000;
12'b010010101010: dataB <= 32'b00000010111101000100100101011010;
12'b010010101011: dataB <= 32'b00000110011110000010101000101101;
12'b010010101100: dataB <= 32'b01001111101101100101010010001101;
12'b010010101101: dataB <= 32'b00001001000011110001010101001101;
12'b010010101110: dataB <= 32'b10100100111011110011111101101101;
12'b010010101111: dataB <= 32'b00000101100111011010110010000010;
12'b010010110000: dataB <= 32'b00110001000011010100011001000100;
12'b010010110001: dataB <= 32'b00000001001100001011000111100110;
12'b010010110010: dataB <= 32'b00000000000010101110011000110101;
12'b010010110011: dataB <= 32'b00000000000000000000000000000000;
12'b010010110100: dataB <= 32'b01101011101111101101101101011011;
12'b010010110101: dataB <= 32'b00000111101001100101011001101000;
12'b010010110110: dataB <= 32'b10001101101110111001001100001001;
12'b010010110111: dataB <= 32'b00000010000101000110110001010110;
12'b010010111000: dataB <= 32'b00111101000100111011010011110010;
12'b010010111001: dataB <= 32'b00000100100010010110101111110011;
12'b010010111010: dataB <= 32'b01101001010111010011111010110001;
12'b010010111011: dataB <= 32'b00000101010011010101100110001000;
12'b010010111100: dataB <= 32'b11010111111001011010100101101111;
12'b010010111101: dataB <= 32'b00001011110100110001110000111001;
12'b010010111110: dataB <= 32'b11100101000001111000011000101000;
12'b010010111111: dataB <= 32'b00000110001001100001111010010010;
12'b010011000000: dataB <= 32'b01011011001000111100000010010101;
12'b010011000001: dataB <= 32'b00000111011001001110100101101011;
12'b010011000010: dataB <= 32'b10101110011000101100110010111001;
12'b010011000011: dataB <= 32'b00000011000100010111010011110010;
12'b010011000100: dataB <= 32'b11100100011110100001101000101100;
12'b010011000101: dataB <= 32'b00001010111110011010100111011100;
12'b010011000110: dataB <= 32'b11000101000000010010000010111010;
12'b010011000111: dataB <= 32'b00000101001010001010010000011010;
12'b010011001000: dataB <= 32'b01101011100000111011010000101111;
12'b010011001001: dataB <= 32'b00000101001100010111100011011110;
12'b010011001010: dataB <= 32'b00101011000110000100000110101010;
12'b010011001011: dataB <= 32'b00000100000011011111110110100011;
12'b010011001100: dataB <= 32'b00011011111010111000101001000001;
12'b010011001101: dataB <= 32'b00000101101101010010100001000011;
12'b010011001110: dataB <= 32'b10110011010101111101100101101010;
12'b010011001111: dataB <= 32'b00000101111110001011101011110100;
12'b010011010000: dataB <= 32'b11101100110101110001111001011100;
12'b010011010001: dataB <= 32'b00000111000001100011000011001100;
12'b010011010010: dataB <= 32'b00111101000010100000011010000111;
12'b010011010011: dataB <= 32'b00001001100011101000101111010001;
12'b010011010100: dataB <= 32'b10110111101011101101101000001001;
12'b010011010101: dataB <= 32'b00000011001001001110111011000010;
12'b010011010110: dataB <= 32'b00101000101110011100011000101100;
12'b010011010111: dataB <= 32'b00001100110101100111000111010011;
12'b010011011000: dataB <= 32'b10001000111001000000100110111001;
12'b010011011001: dataB <= 32'b00001111010001101110111000111100;
12'b010011011010: dataB <= 32'b11011011100101001000100111010000;
12'b010011011011: dataB <= 32'b00001010000001110001001101010011;
12'b010011011100: dataB <= 32'b01100111011100111100100101011101;
12'b010011011101: dataB <= 32'b00001100001100101111000110001100;
12'b010011011110: dataB <= 32'b01100110100110010000011000001000;
12'b010011011111: dataB <= 32'b00000111100111100011001110111001;
12'b010011100000: dataB <= 32'b01100010101011001101101000100100;
12'b010011100001: dataB <= 32'b00000010101001001001011111000101;
12'b010011100010: dataB <= 32'b11000010111000110001000011101100;
12'b010011100011: dataB <= 32'b00000111100101100111100101011100;
12'b010011100100: dataB <= 32'b10100110110110001101011000111101;
12'b010011100101: dataB <= 32'b00000111010101011011101110111010;
12'b010011100110: dataB <= 32'b11101100110101000101110000101011;
12'b010011100111: dataB <= 32'b00001010001000110011010110101001;
12'b010011101000: dataB <= 32'b00110111000110000001101000001011;
12'b010011101001: dataB <= 32'b00000100001011010111011011101010;
12'b010011101010: dataB <= 32'b11001011001101011110100100011100;
12'b010011101011: dataB <= 32'b00001100000101101011000100111101;
12'b010011101100: dataB <= 32'b01010100100000011010000011110100;
12'b010011101101: dataB <= 32'b00001001001101100101001010001111;
12'b010011101110: dataB <= 32'b11101101000101001010000110111100;
12'b010011101111: dataB <= 32'b00000100101100000100101010010000;
12'b010011110000: dataB <= 32'b11010011000101101100100111011000;
12'b010011110001: dataB <= 32'b00000110011110010011110101000010;
12'b010011110010: dataB <= 32'b10011110101000101010000000101101;
12'b010011110011: dataB <= 32'b00001110011000100000111111000110;
12'b010011110100: dataB <= 32'b01100011100101001011110100010101;
12'b010011110101: dataB <= 32'b00000101111011000111001001100000;
12'b010011110110: dataB <= 32'b10010001101001101110000100111100;
12'b010011110111: dataB <= 32'b00001011001000101011010001100111;
12'b010011111000: dataB <= 32'b10001000101010101011111011111011;
12'b010011111001: dataB <= 32'b00001010110111011110110101011011;
12'b010011111010: dataB <= 32'b10011011111010111000101101111001;
12'b010011111011: dataB <= 32'b00001000001000100010110101011101;
12'b010011111100: dataB <= 32'b11100101110001010010000111111001;
12'b010011111101: dataB <= 32'b00000101101101011111011101101010;
12'b010011111110: dataB <= 32'b01100111000011100110001100010110;
12'b010011111111: dataB <= 32'b00001110001000110100110110010000;
12'b010100000000: dataB <= 32'b10000010110101000100010100011000;
12'b010100000001: dataB <= 32'b00000101011101000110100000101100;
12'b010100000010: dataB <= 32'b00001011100101011101000010101010;
12'b010100000011: dataB <= 32'b00001010000100101111011101000101;
12'b010100000100: dataB <= 32'b10100100111111110100101101101111;
12'b010100000101: dataB <= 32'b00000110100110011010110010001010;
12'b010100000110: dataB <= 32'b10101111000111010100111010100101;
12'b010100000111: dataB <= 32'b00000001101010001010111111010110;
12'b010100001000: dataB <= 32'b00000000000010011110101000010110;
12'b010100001001: dataB <= 32'b00000000000000000000000000000000;
12'b010100001010: dataB <= 32'b01100111110011100110001011111100;
12'b010100001011: dataB <= 32'b00001000001001100011011010000000;
12'b010100001100: dataB <= 32'b01001001100111010001011100101011;
12'b010100001101: dataB <= 32'b00000011100011001000101001000110;
12'b010100001110: dataB <= 32'b11111101010001000010110011110000;
12'b010100001111: dataB <= 32'b00000110000001011000101011110011;
12'b010100010000: dataB <= 32'b01100111011011010100101010110010;
12'b010100010001: dataB <= 32'b00000101010010010001011110100000;
12'b010100010010: dataB <= 32'b01010001110101100010010101101110;
12'b010100010011: dataB <= 32'b00001011010110101101110101000001;
12'b010100010100: dataB <= 32'b11100101000010010000011001101000;
12'b010100010101: dataB <= 32'b00000110101001011011111010011010;
12'b010100010110: dataB <= 32'b01011011001000111011100001110011;
12'b010100010111: dataB <= 32'b00000110011001010010011101101011;
12'b010100011000: dataB <= 32'b01110010100000101100010001110111;
12'b010100011001: dataB <= 32'b00000100100010010101001111110011;
12'b010100011010: dataB <= 32'b01101000100010110001111001001100;
12'b010100011011: dataB <= 32'b00001001011110011100100111010101;
12'b010100011100: dataB <= 32'b01000100111000100001100001111000;
12'b010100011101: dataB <= 32'b00000101101001010000001100100010;
12'b010100011110: dataB <= 32'b11100111100101000010110000101100;
12'b010100011111: dataB <= 32'b00000101101011010011011111001110;
12'b010100100000: dataB <= 32'b01101011001010000100000111001010;
12'b010100100001: dataB <= 32'b00000101000001011011110110100011;
12'b010100100010: dataB <= 32'b11010101110111001001001010000001;
12'b010100100011: dataB <= 32'b00000110001100010110011101001010;
12'b010100100100: dataB <= 32'b00101111011101110101100110001001;
12'b010100100101: dataB <= 32'b00000100011100000111100011110101;
12'b010100100110: dataB <= 32'b01101100111010000001101000011101;
12'b010100100111: dataB <= 32'b00001000100001100011000011000101;
12'b010100101000: dataB <= 32'b11111101001110111000101011001000;
12'b010100101001: dataB <= 32'b00001010100100101010110011100001;
12'b010100101010: dataB <= 32'b00110001110011100110001000101001;
12'b010100101011: dataB <= 32'b00000100000111001110110011001011;
12'b010100101100: dataB <= 32'b10101010110010011100011000101100;
12'b010100101101: dataB <= 32'b00001100010111100111001011010011;
12'b010100101110: dataB <= 32'b00001010110001011000010101111000;
12'b010100101111: dataB <= 32'b00001111010100110001000000111100;
12'b010100110000: dataB <= 32'b10010111100001100000010111010000;
12'b010100110001: dataB <= 32'b00001011100010101111010101010011;
12'b010100110010: dataB <= 32'b01100011011100111100000100011011;
12'b010100110011: dataB <= 32'b00001100001110101111001110001100;
12'b010100110100: dataB <= 32'b11101000101010100000011001001000;
12'b010100110101: dataB <= 32'b00001000100111100001001111001001;
12'b010100110110: dataB <= 32'b11100100101010111110001001100100;
12'b010100110111: dataB <= 32'b00000011100111000111010110110101;
12'b010100111000: dataB <= 32'b10000100101101001000100100001010;
12'b010100111001: dataB <= 32'b00001001000101100011100101011100;
12'b010100111010: dataB <= 32'b00100110111010000101010111111101;
12'b010100111011: dataB <= 32'b00000110110101010111101011000011;
12'b010100111100: dataB <= 32'b01101100111000111101010001001000;
12'b010100111101: dataB <= 32'b00001011001001101111011110111010;
12'b010100111110: dataB <= 32'b11110101001110010001101000101011;
12'b010100111111: dataB <= 32'b00000100101001010101010111110010;
12'b010101000000: dataB <= 32'b01001011000101001110010010111010;
12'b010101000001: dataB <= 32'b00001101000110101011001000110101;
12'b010101000010: dataB <= 32'b01011000011100100001100011010010;
12'b010101000011: dataB <= 32'b00001001001101100101001001111111;
12'b010101000100: dataB <= 32'b00101101001001011001110101111011;
12'b010101000101: dataB <= 32'b00000101001011000110011110100001;
12'b010101000110: dataB <= 32'b01010000111101101100100110011000;
12'b010101000111: dataB <= 32'b00000100111101001111110001001010;
12'b010101001000: dataB <= 32'b00100000101000111001100001001010;
12'b010101001001: dataB <= 32'b00001101011010100000111110110111;
12'b010101001010: dataB <= 32'b01011111101001001011100011110011;
12'b010101001011: dataB <= 32'b00000100111010000101000001111000;
12'b010101001100: dataB <= 32'b01001101100001011101110011111010;
12'b010101001101: dataB <= 32'b00001011101010101001010101001111;
12'b010101001110: dataB <= 32'b01001100011110101100001010111100;
12'b010101001111: dataB <= 32'b00001001111000011110110101011011;
12'b010101010000: dataB <= 32'b01010101110111001001001100111011;
12'b010101010001: dataB <= 32'b00001001001000100010110101010101;
12'b010101010010: dataB <= 32'b11100001110101100001110110111001;
12'b010101010011: dataB <= 32'b00000110001100011011011101110010;
12'b010101010100: dataB <= 32'b01100111000011010110101011011000;
12'b010101010101: dataB <= 32'b00001111001010110110111110100000;
12'b010101010110: dataB <= 32'b00000100101000111011110011010110;
12'b010101010111: dataB <= 32'b00000011111100001010010100100100;
12'b010101011000: dataB <= 32'b10000111011101010100110011001000;
12'b010101011001: dataB <= 32'b00001011000101101011100001000100;
12'b010101011010: dataB <= 32'b10100100111111101101011101110001;
12'b010101011011: dataB <= 32'b00000111100110011100110010010010;
12'b010101011100: dataB <= 32'b00101111001111001101011011100110;
12'b010101011101: dataB <= 32'b00000010101000001010110011000111;
12'b010101011110: dataB <= 32'b00000000000010001110100111110110;
12'b010101011111: dataB <= 32'b00000000000000000000000000000000;
12'b010101100000: dataB <= 32'b11111000110011000000111110001000;
12'b010101100001: dataB <= 32'b00000100101111101100111000001011;
12'b010101100010: dataB <= 32'b11110011101100101001010101100110;
12'b010101100011: dataB <= 32'b00000001111000010101101111001101;
12'b010101100100: dataB <= 32'b01101000000101011101111000011000;
12'b010101100101: dataB <= 32'b00000000110011010101001101111000;
12'b010101100110: dataB <= 32'b11101100110010010001011001001010;
12'b010101100111: dataB <= 32'b00001001010101101111011100001010;
12'b010101101000: dataB <= 32'b11111011011101001100110111010100;
12'b010101101001: dataB <= 32'b00001011001001111010100100101101;
12'b010101101010: dataB <= 32'b00100000110100001011010100001100;
12'b010101101011: dataB <= 32'b00000100110010111101001001011011;
12'b010101101100: dataB <= 32'b10100101001001110110001001111100;
12'b010101101101: dataB <= 32'b00001100110011001111011001101100;
12'b010101101110: dataB <= 32'b01010000011010001110101011111100;
12'b010101101111: dataB <= 32'b00000001010110100111010101101000;
12'b010101110000: dataB <= 32'b01010000101100111010010110001101;
12'b010101110001: dataB <= 32'b00001111001101010011000110101001;
12'b010101110010: dataB <= 32'b11011101110100110110111100011100;
12'b010101110011: dataB <= 32'b00000100110100000111011101001110;
12'b010101110100: dataB <= 32'b10110010110001011101110110011110;
12'b010101110101: dataB <= 32'b00000101110100101111011011011001;
12'b010101110110: dataB <= 32'b11100100101010000011110101010001;
12'b010101110111: dataB <= 32'b00000000110101111011001001101010;
12'b010101111000: dataB <= 32'b10111011010100100001100000101011;
12'b010101111001: dataB <= 32'b00000110010011001111010001011101;
12'b010101111010: dataB <= 32'b01101110100010110100010100110011;
12'b010101111011: dataB <= 32'b00001110010111110001110010100000;
12'b010101111100: dataB <= 32'b11011100100100110011111110101111;
12'b010101111101: dataB <= 32'b00000000101110100000111010101001;
12'b010101111110: dataB <= 32'b11100110000100010010000100001001;
12'b010101111111: dataB <= 32'b00000010001010011000101000111000;
12'b010110000000: dataB <= 32'b10111000011111000000110100101110;
12'b010110000001: dataB <= 32'b00000011110111011001100001100001;
12'b010110000010: dataB <= 32'b01011000101010001011000110001110;
12'b010110000011: dataB <= 32'b00001011100111100100110001110001;
12'b010110000100: dataB <= 32'b00011001101000001101001100010100;
12'b010110000101: dataB <= 32'b00001010000001100000011110000110;
12'b010110000110: dataB <= 32'b01110001010000001100111000010001;
12'b010110000111: dataB <= 32'b00000001001000101010100001110101;
12'b010110001000: dataB <= 32'b10101110111010000110001101110111;
12'b010110001001: dataB <= 32'b00000111000111100110100010001011;
12'b010110001010: dataB <= 32'b10010100101100001010110100001101;
12'b010110001011: dataB <= 32'b00000011101110100110111100111001;
12'b010110001100: dataB <= 32'b01010100110111000010000010001100;
12'b010110001101: dataB <= 32'b00000011111000101011110010111010;
12'b010110001110: dataB <= 32'b00010111110100010101100101010111;
12'b010110001111: dataB <= 32'b00000010101101110010111010010101;
12'b010110010000: dataB <= 32'b11011100110010101011111110110000;
12'b010110010001: dataB <= 32'b00001010110010110101010001100001;
12'b010110010010: dataB <= 32'b00011100100110101110000100011101;
12'b010110010011: dataB <= 32'b00000100101001101110100001001010;
12'b010110010100: dataB <= 32'b01100110010100110011010101101110;
12'b010110010101: dataB <= 32'b00000100110110101011010101011000;
12'b010110010110: dataB <= 32'b01100011101011001101101101011010;
12'b010110010111: dataB <= 32'b00000011000101100100101010101110;
12'b010110011000: dataB <= 32'b00001111001100110110111001011001;
12'b010110011001: dataB <= 32'b00000110101101100100110111101100;
12'b010110011010: dataB <= 32'b11100100100100111101001101110100;
12'b010110011011: dataB <= 32'b00000101110101001111110000100010;
12'b010110011100: dataB <= 32'b10011111011110010100101100010011;
12'b010110011101: dataB <= 32'b00001110110110111001100001001101;
12'b010110011110: dataB <= 32'b01010100111100110110000101011101;
12'b010110011111: dataB <= 32'b00001101000101011110111111100010;
12'b010110100000: dataB <= 32'b00110101000001110101101001111000;
12'b010110100001: dataB <= 32'b00001101010110100001110100001100;
12'b010110100010: dataB <= 32'b10110001100110111101001101011000;
12'b010110100011: dataB <= 32'b00000101001000101010101111101101;
12'b010110100100: dataB <= 32'b00001111100110000010101110001010;
12'b010110100101: dataB <= 32'b00001100001100011011000001101101;
12'b010110100110: dataB <= 32'b01111011010100100001101101100110;
12'b010110100111: dataB <= 32'b00000100001101011010111010101101;
12'b010110101000: dataB <= 32'b01111010111100111100111100110010;
12'b010110101001: dataB <= 32'b00000110010011101111001001011100;
12'b010110101010: dataB <= 32'b11100000110011010001011100001001;
12'b010110101011: dataB <= 32'b00000101000001011110010000001010;
12'b010110101100: dataB <= 32'b11010101110101111110001011011001;
12'b010110101101: dataB <= 32'b00001110011000001011101010000110;
12'b010110101110: dataB <= 32'b11101111110010011101010100011001;
12'b010110101111: dataB <= 32'b00000010101001110000101010010101;
12'b010110110000: dataB <= 32'b01011110110110101000101000100100;
12'b010110110001: dataB <= 32'b00000011010000011001000101010011;
12'b010110110010: dataB <= 32'b11100110100010101001100011001000;
12'b010110110011: dataB <= 32'b00000100011010011001101011100001;
12'b010110110100: dataB <= 32'b00000000000011010011101011010000;
12'b010110110101: dataB <= 32'b00000000000000000000000000000000;
12'b010110110110: dataB <= 32'b10110110101010110000101101100101;
12'b010110110111: dataB <= 32'b00000100110000101100110100001100;
12'b010110111000: dataB <= 32'b01110111100100100010000100100111;
12'b010110111001: dataB <= 32'b00000010111011011001110011010101;
12'b010110111010: dataB <= 32'b01100010000101101110001001011000;
12'b010110111011: dataB <= 32'b00000001010110010111010001100000;
12'b010110111100: dataB <= 32'b10101010101101111001011000101010;
12'b010110111101: dataB <= 32'b00001001110101110011010100001011;
12'b010110111110: dataB <= 32'b00111101010001010101000111110100;
12'b010110111111: dataB <= 32'b00001010001000111000011100111110;
12'b010111000000: dataB <= 32'b01100000110100001100000100001110;
12'b010111000001: dataB <= 32'b00000100110011111100111101011011;
12'b010111000010: dataB <= 32'b10100101001010000110001010111011;
12'b010111000011: dataB <= 32'b00001100110001010011100001101100;
12'b010111000100: dataB <= 32'b01001100100010011110101100111010;
12'b010111000101: dataB <= 32'b00000010011001101001010001010000;
12'b010111000110: dataB <= 32'b00001110110100110010110110001110;
12'b010111000111: dataB <= 32'b00001111001010010011001010011001;
12'b010111001000: dataB <= 32'b00100001110101000111011101011010;
12'b010111001001: dataB <= 32'b00000101010101001001101001011111;
12'b010111001010: dataB <= 32'b00110000101001101110000111111110;
12'b010111001011: dataB <= 32'b00000110010101110001010011001001;
12'b010111001100: dataB <= 32'b11100010101010000011110101010010;
12'b010111001101: dataB <= 32'b00000001110111111011000001100010;
12'b010111001110: dataB <= 32'b11111101001000010010000000101101;
12'b010111001111: dataB <= 32'b00000110110100010001011001100101;
12'b010111010000: dataB <= 32'b01101010011010110100000101010100;
12'b010111010001: dataB <= 32'b00001111010100110101101010010000;
12'b010111010010: dataB <= 32'b10011010100100111100011110001101;
12'b010111010011: dataB <= 32'b00000000110001100000111010011001;
12'b010111010100: dataB <= 32'b01100000000100001010110011101011;
12'b010111010101: dataB <= 32'b00000001101100010110101100100001;
12'b010111010110: dataB <= 32'b11110100010010110000100100101111;
12'b010111010111: dataB <= 32'b00000100111001011101100001010001;
12'b010111011000: dataB <= 32'b01010110101110001011000110001110;
12'b010111011001: dataB <= 32'b00001010100110100010110001100001;
12'b010111011010: dataB <= 32'b00011101101100010101111100110010;
12'b010111011011: dataB <= 32'b00001000100001011100100010010110;
12'b010111011100: dataB <= 32'b01110011001000010101101000010001;
12'b010111011101: dataB <= 32'b00000000101011100110011101111101;
12'b010111011110: dataB <= 32'b10101110110010010110001110110101;
12'b010111011111: dataB <= 32'b00000110000111100010100010001011;
12'b010111100000: dataB <= 32'b00010010110000001011010100001111;
12'b010111100001: dataB <= 32'b00000011110000100110111000101010;
12'b010111100010: dataB <= 32'b11010100111010110001100010001110;
12'b010111100011: dataB <= 32'b00000100111010101111101110101001;
12'b010111100100: dataB <= 32'b00011101111000100110010110011000;
12'b010111100101: dataB <= 32'b00000010110000110010110010011101;
12'b010111100110: dataB <= 32'b00011010110010101011101110101110;
12'b010111100111: dataB <= 32'b00001010110001110111001001010010;
12'b010111101000: dataB <= 32'b10011010100110111101110101111110;
12'b010111101001: dataB <= 32'b00000100001011101010011000111010;
12'b010111101010: dataB <= 32'b10100010010000110011110101101111;
12'b010111101011: dataB <= 32'b00000101110111101101010001000000;
12'b010111101100: dataB <= 32'b00100111101011010101001110010111;
12'b010111101101: dataB <= 32'b00000010100111100010101010111110;
12'b010111101110: dataB <= 32'b10010001010101000111001010011000;
12'b010111101111: dataB <= 32'b00000110101101100100110111101011;
12'b010111110000: dataB <= 32'b01100010100101000101101110010010;
12'b010111110001: dataB <= 32'b00000110010110010101110100011011;
12'b010111110010: dataB <= 32'b11100011011010010100101100010001;
12'b010111110011: dataB <= 32'b00001111010011111011011001011101;
12'b010111110100: dataB <= 32'b11010101000001000110100110111110;
12'b010111110101: dataB <= 32'b00001100000011011110111111010001;
12'b010111110110: dataB <= 32'b11110010111001111101101010110111;
12'b010111110111: dataB <= 32'b00001101110100100101110000001100;
12'b010111111000: dataB <= 32'b11110101011111000100101110010110;
12'b010111111001: dataB <= 32'b00000100001001101000101011110100;
12'b010111111010: dataB <= 32'b00010101101101111010101101101000;
12'b010111111011: dataB <= 32'b00001011101010011011000001110101;
12'b010111111100: dataB <= 32'b00111101001000010010001100100100;
12'b010111111101: dataB <= 32'b00000100001111011010111010110101;
12'b010111111110: dataB <= 32'b10111000110101000101011100110000;
12'b010111111111: dataB <= 32'b00000110110100101111000001011100;
12'b011000000000: dataB <= 32'b01100000110011000000111011000111;
12'b011000000001: dataB <= 32'b00000100000011011010010100001011;
12'b011000000010: dataB <= 32'b10011011111010001101111100010111;
12'b011000000011: dataB <= 32'b00001110110101010001110010010110;
12'b011000000100: dataB <= 32'b11110011101010100101000101011010;
12'b011000000101: dataB <= 32'b00000010001011101110100010100101;
12'b011000000110: dataB <= 32'b10011110110110010000010111100100;
12'b011000000111: dataB <= 32'b00000011010010011001001001010011;
12'b011000001000: dataB <= 32'b01100010100010011001010010101010;
12'b011000001001: dataB <= 32'b00000101011100011111101011010001;
12'b011000001010: dataB <= 32'b00000000000011010011001011001111;
12'b011000001011: dataB <= 32'b00000000000000000000000000000000;
12'b011000001100: dataB <= 32'b01110100100010011000011100000011;
12'b011000001101: dataB <= 32'b00000101010001101010101100001101;
12'b011000001110: dataB <= 32'b10111001011100010010100011101001;
12'b011000001111: dataB <= 32'b00000100011100011111110111011100;
12'b011000010000: dataB <= 32'b10011100000101110110001010010111;
12'b011000010001: dataB <= 32'b00000001111000011001010101001000;
12'b011000010010: dataB <= 32'b01101000101001101001011000001010;
12'b011000010011: dataB <= 32'b00001010010100110011001100001100;
12'b011000010100: dataB <= 32'b10111101000101011101011000010100;
12'b011000010101: dataB <= 32'b00001001100111110100010101001110;
12'b011000010110: dataB <= 32'b10011110110100001100110011101111;
12'b011000010111: dataB <= 32'b00000101010101111100110001010011;
12'b011000011000: dataB <= 32'b11100111000110010101111011111010;
12'b011000011001: dataB <= 32'b00001100101111010101100101110100;
12'b011000011010: dataB <= 32'b11001010101010101110011101111000;
12'b011000011011: dataB <= 32'b00000011011011101011001101000000;
12'b011000011100: dataB <= 32'b11001110111000101011010101101110;
12'b011000011101: dataB <= 32'b00001110001000010101010010001000;
12'b011000011110: dataB <= 32'b01100111110001011111101110011000;
12'b011000011111: dataB <= 32'b00000101110110001111110001110111;
12'b011000100000: dataB <= 32'b11101110100001110110001001011110;
12'b011000100001: dataB <= 32'b00000110110101110011001010111000;
12'b011000100010: dataB <= 32'b00100000101010000011110101110011;
12'b011000100011: dataB <= 32'b00000010111010111010110101011011;
12'b011000100100: dataB <= 32'b11111101000000001010110000110000;
12'b011000100101: dataB <= 32'b00000110110100010011011101110101;
12'b011000100110: dataB <= 32'b01100110011010110011100101110101;
12'b011000100111: dataB <= 32'b00001111010010111001100001111000;
12'b011000101000: dataB <= 32'b10010110101000111100111101101010;
12'b011000101001: dataB <= 32'b00000000110100100000111010001001;
12'b011000101010: dataB <= 32'b00011010000100001011100011001101;
12'b011000101011: dataB <= 32'b00000001001111010100110000011010;
12'b011000101100: dataB <= 32'b00101110001110011000010100110001;
12'b011000101101: dataB <= 32'b00000101111010100001100001000010;
12'b011000101110: dataB <= 32'b10010100110010000011000110001111;
12'b011000101111: dataB <= 32'b00001001100101100010101101010001;
12'b011000110000: dataB <= 32'b11100001101100100110011100110000;
12'b011000110001: dataB <= 32'b00000111000001011010100010100101;
12'b011000110010: dataB <= 32'b01110011000000011110001000010001;
12'b011000110011: dataB <= 32'b00000000101110100010011010000101;
12'b011000110100: dataB <= 32'b10101100101110100101111110110010;
12'b011000110101: dataB <= 32'b00000101001000100000011110001011;
12'b011000110110: dataB <= 32'b10010010110100001100000100010000;
12'b011000110111: dataB <= 32'b00000100010010100110111000100010;
12'b011000111000: dataB <= 32'b10010100111110100001010001110000;
12'b011000111001: dataB <= 32'b00000101111011110011100110100001;
12'b011000111010: dataB <= 32'b11100001111000110110110111011001;
12'b011000111011: dataB <= 32'b00000010110010110000101010100100;
12'b011000111100: dataB <= 32'b01011010110010101011011110001011;
12'b011000111101: dataB <= 32'b00001010110000110111000001001010;
12'b011000111110: dataB <= 32'b11010110101011000101010111011110;
12'b011000111111: dataB <= 32'b00000011101100100110011000110010;
12'b011001000000: dataB <= 32'b00011110010000110100010101110000;
12'b011001000001: dataB <= 32'b00000110011000101111001000110001;
12'b011001000010: dataB <= 32'b10101011100111011100011111010101;
12'b011001000011: dataB <= 32'b00000001101010100000101011001101;
12'b011001000100: dataB <= 32'b11010011011001011111101011010111;
12'b011001000101: dataB <= 32'b00000110001110100010110011100010;
12'b011001000110: dataB <= 32'b11011110100101001101111110010000;
12'b011001000111: dataB <= 32'b00000110110110011001111000011011;
12'b011001001000: dataB <= 32'b00100101011010011100011100001111;
12'b011001001001: dataB <= 32'b00001111010000111101001101100110;
12'b011001001010: dataB <= 32'b01010111000101010110110111111110;
12'b011001001011: dataB <= 32'b00001011000010011110111111001001;
12'b011001001100: dataB <= 32'b10110010110010001101101011010110;
12'b011001001101: dataB <= 32'b00001110010010101011101100010101;
12'b011001001110: dataB <= 32'b00110111010111000100011110110100;
12'b011001001111: dataB <= 32'b00000011101011100110100111110100;
12'b011001010000: dataB <= 32'b00011001110001110010111100100110;
12'b011001010001: dataB <= 32'b00001011001001011011000101111101;
12'b011001010010: dataB <= 32'b10111100111100001010111011100011;
12'b011001010011: dataB <= 32'b00000100010000011010111110111100;
12'b011001010100: dataB <= 32'b11110110101001001101101100101110;
12'b011001010101: dataB <= 32'b00000110110100101110111101100100;
12'b011001010110: dataB <= 32'b00011110110010101000101010100110;
12'b011001010111: dataB <= 32'b00000010100101010110010100001100;
12'b011001011000: dataB <= 32'b10011111111010010101111101010101;
12'b011001011001: dataB <= 32'b00001111010011010101111010100110;
12'b011001011010: dataB <= 32'b10110111100010101100110110111011;
12'b011001011011: dataB <= 32'b00000001101101101010011110101101;
12'b011001011100: dataB <= 32'b11011100110101111000010110100100;
12'b011001011101: dataB <= 32'b00000011110100011001001001010011;
12'b011001011110: dataB <= 32'b11100000011110001001010010001101;
12'b011001011111: dataB <= 32'b00000110011101100011101011000000;
12'b011001100000: dataB <= 32'b00000000000011001010101010101110;
12'b011001100001: dataB <= 32'b00000000000000000000000000000000;
12'b011001100010: dataB <= 32'b11110000011010000000011011000010;
12'b011001100011: dataB <= 32'b00000101010011101000101000011101;
12'b011001100100: dataB <= 32'b00111101010000010011010011001010;
12'b011001100101: dataB <= 32'b00000101011110100011110011100100;
12'b011001100110: dataB <= 32'b11010110000110000110001010110110;
12'b011001100111: dataB <= 32'b00000010111010011011011000111000;
12'b011001101000: dataB <= 32'b00100110100101011001100111101010;
12'b011001101001: dataB <= 32'b00001010110011110101000100001101;
12'b011001101010: dataB <= 32'b11111100111001100101101000010100;
12'b011001101011: dataB <= 32'b00001000100110101110001101011110;
12'b011001101100: dataB <= 32'b11011110110100010101100100010001;
12'b011001101101: dataB <= 32'b00000101110101111010100101010011;
12'b011001101110: dataB <= 32'b11100111000110011101111100111000;
12'b011001101111: dataB <= 32'b00001100101101011001101001110100;
12'b011001110000: dataB <= 32'b01001000110010110110001110010110;
12'b011001110001: dataB <= 32'b00000100011101101101001000101001;
12'b011001110010: dataB <= 32'b11001111000000101011110101101111;
12'b011001110011: dataB <= 32'b00001101000101010111010101111000;
12'b011001110100: dataB <= 32'b01101011101101110111101110110101;
12'b011001110101: dataB <= 32'b00000110110111010011110110000111;
12'b011001110110: dataB <= 32'b01101010011110000110001010111110;
12'b011001110111: dataB <= 32'b00000111010110110011000010100000;
12'b011001111000: dataB <= 32'b01011110101010000011110101110100;
12'b011001111001: dataB <= 32'b00000011111100111000101001011011;
12'b011001111010: dataB <= 32'b11111100110100001011100000110011;
12'b011001111011: dataB <= 32'b00000111010100010111100001111101;
12'b011001111100: dataB <= 32'b01100010010110101011010110010110;
12'b011001111101: dataB <= 32'b00001111001111111011010101100000;
12'b011001111110: dataB <= 32'b10010100101101000101001101001000;
12'b011001111111: dataB <= 32'b00000001010111100000111001111001;
12'b011010000000: dataB <= 32'b10010100000100001100010011001111;
12'b011010000001: dataB <= 32'b00000001110001010010110100001010;
12'b011010000010: dataB <= 32'b10101010000110000000010101010010;
12'b011010000011: dataB <= 32'b00000110111011100011100000111010;
12'b011010000100: dataB <= 32'b11010010110101111011000110010000;
12'b011010000101: dataB <= 32'b00001000100100100000101101001001;
12'b011010000110: dataB <= 32'b10100101101000110110111100101110;
12'b011010000111: dataB <= 32'b00000101100001010110100110101101;
12'b011010001000: dataB <= 32'b01110010111000101110101000110001;
12'b011010001001: dataB <= 32'b00000000110001100000011010001101;
12'b011010001010: dataB <= 32'b01101010101010101101101111001111;
12'b011010001011: dataB <= 32'b00000100101001011100100010000011;
12'b011010001100: dataB <= 32'b01010000111100001100110100010010;
12'b011010001101: dataB <= 32'b00000100010011100110110100011011;
12'b011010001110: dataB <= 32'b10010101000010010001000010010011;
12'b011010001111: dataB <= 32'b00000111011011110111011110010001;
12'b011010010000: dataB <= 32'b10100111110101000111010111111001;
12'b011010010001: dataB <= 32'b00000011010100101110100010100100;
12'b011010010010: dataB <= 32'b10011000110110100011001101101001;
12'b011010010011: dataB <= 32'b00001010101111110110111000111010;
12'b011010010100: dataB <= 32'b01010100101111001100111000111110;
12'b011010010101: dataB <= 32'b00000011001110100010010100110011;
12'b011010010110: dataB <= 32'b10011010010100111100110101110000;
12'b011010010111: dataB <= 32'b00000111011001101111000100100001;
12'b011010011000: dataB <= 32'b00101101100011011011111111010010;
12'b011010011001: dataB <= 32'b00000001001100011110101011010101;
12'b011010011010: dataB <= 32'b01010101100001101111101011110110;
12'b011010011011: dataB <= 32'b00000110001110100010110011011010;
12'b011010011100: dataB <= 32'b10011100100101011110001110001101;
12'b011010011101: dataB <= 32'b00000111110111011111111000011100;
12'b011010011110: dataB <= 32'b01100111011010011100011100001110;
12'b011010011111: dataB <= 32'b00001111001101111101000001110110;
12'b011010100000: dataB <= 32'b11010111001001101111001001011110;
12'b011010100001: dataB <= 32'b00001001100001011110111110110000;
12'b011010100010: dataB <= 32'b00110000101010010101011100010101;
12'b011010100011: dataB <= 32'b00001110001111101111101000011110;
12'b011010100100: dataB <= 32'b01111001001011000011111111010001;
12'b011010100101: dataB <= 32'b00000011101100100100100111110011;
12'b011010100110: dataB <= 32'b00011101110001101010111011100100;
12'b011010100111: dataB <= 32'b00001010100111011011000110000101;
12'b011010101000: dataB <= 32'b01111100110100001011101010000001;
12'b011010101001: dataB <= 32'b00000100010010011010111110111100;
12'b011010101010: dataB <= 32'b11110100100001010110001100001100;
12'b011010101011: dataB <= 32'b00000111010100101110110101100100;
12'b011010101100: dataB <= 32'b11011100110110010000011001100101;
12'b011010101101: dataB <= 32'b00000001100111010010011000001100;
12'b011010101110: dataB <= 32'b01100101111010100101101101010011;
12'b011010101111: dataB <= 32'b00001111010000011011111010110110;
12'b011010110000: dataB <= 32'b00111001011010110100100111111100;
12'b011010110001: dataB <= 32'b00000001110000100110011010110101;
12'b011010110010: dataB <= 32'b00011100110101101000010101100101;
12'b011010110011: dataB <= 32'b00000100010110011011001101010100;
12'b011010110100: dataB <= 32'b10011100100001110001010001101111;
12'b011010110101: dataB <= 32'b00000111111101100111101010101000;
12'b011010110110: dataB <= 32'b00000000000011000010011010101100;
12'b011010110111: dataB <= 32'b00000000000000000000000000000000;
12'b011010111000: dataB <= 32'b10101100010001101000011001100001;
12'b011010111001: dataB <= 32'b00000101110100100110100100101110;
12'b011010111010: dataB <= 32'b10111101001000001011110010101100;
12'b011010111011: dataB <= 32'b00000110111110101001110011011011;
12'b011010111100: dataB <= 32'b01010000001010010110001011010101;
12'b011010111101: dataB <= 32'b00000100011100011101011000101001;
12'b011010111110: dataB <= 32'b11100100100001010001110111001010;
12'b011010111111: dataB <= 32'b00001010110010110100111100010101;
12'b011011000000: dataB <= 32'b00111100101101101101111000110100;
12'b011011000001: dataB <= 32'b00000111100110101010000101101111;
12'b011011000010: dataB <= 32'b00011110110100011110000100010010;
12'b011011000011: dataB <= 32'b00000110110110111000011101010100;
12'b011011000100: dataB <= 32'b11100111000010100101101101110110;
12'b011011000101: dataB <= 32'b00001100001011011101101001111100;
12'b011011000110: dataB <= 32'b11000110111111000101101110110011;
12'b011011000111: dataB <= 32'b00000101111110101101000100011001;
12'b011011001000: dataB <= 32'b00001111001000101100010101110000;
12'b011011001001: dataB <= 32'b00001100000011011001011001100001;
12'b011011001010: dataB <= 32'b01110001101010001111101111010010;
12'b011011001011: dataB <= 32'b00000111010111011001111010011111;
12'b011011001100: dataB <= 32'b01101000011010010110001011111100;
12'b011011001101: dataB <= 32'b00000111110110110010111110010000;
12'b011011001110: dataB <= 32'b10011100101010000011110110010101;
12'b011011001111: dataB <= 32'b00000100111101110110100001010011;
12'b011011010000: dataB <= 32'b11111010101000001100010001010110;
12'b011011010001: dataB <= 32'b00000111110100011011100110001101;
12'b011011010010: dataB <= 32'b10011110010110101011000110110111;
12'b011011010011: dataB <= 32'b00001111001100111101001001001000;
12'b011011010100: dataB <= 32'b10010010110001001101101100100110;
12'b011011010101: dataB <= 32'b00000010011001011110111001101001;
12'b011011010110: dataB <= 32'b01010000001100001101000011010000;
12'b011011010111: dataB <= 32'b00000001110100010010111000001011;
12'b011011011000: dataB <= 32'b11100100000101101000010101010011;
12'b011011011001: dataB <= 32'b00000111111011100111100000110010;
12'b011011011010: dataB <= 32'b01010010111001110011000110010001;
12'b011011011011: dataB <= 32'b00000111000100011110101100111010;
12'b011011011100: dataB <= 32'b01101001101001000111011100001100;
12'b011011011101: dataB <= 32'b00000100000010010100101010110101;
12'b011011011110: dataB <= 32'b00110000110001000111001000110001;
12'b011011011111: dataB <= 32'b00000000110100011100011010010101;
12'b011011100000: dataB <= 32'b01101000100110110101011110101101;
12'b011011100001: dataB <= 32'b00000100001011011010100010000011;
12'b011011100010: dataB <= 32'b11010001000000010101100100110011;
12'b011011100011: dataB <= 32'b00000100110100100100110000011011;
12'b011011100100: dataB <= 32'b10010101000110000001000010110101;
12'b011011100101: dataB <= 32'b00001000011100111001010110000001;
12'b011011100110: dataB <= 32'b01101101110001011111101000111001;
12'b011011100111: dataB <= 32'b00000011110101101010011110101100;
12'b011011101000: dataB <= 32'b00011000111010011010111100100111;
12'b011011101001: dataB <= 32'b00001010101110110100110000111011;
12'b011011101010: dataB <= 32'b11010010110011010100011010011110;
12'b011011101011: dataB <= 32'b00000011010000011110010100110011;
12'b011011101100: dataB <= 32'b00010110010100111101010101110001;
12'b011011101101: dataB <= 32'b00001000011001101110111100010010;
12'b011011101110: dataB <= 32'b10110001011011011011011111001111;
12'b011011101111: dataB <= 32'b00000001001111011100101011010100;
12'b011011110000: dataB <= 32'b11011001100010000111101100010100;
12'b011011110001: dataB <= 32'b00000110001111100000110011001001;
12'b011011110010: dataB <= 32'b00011010100101101110011101101011;
12'b011011110011: dataB <= 32'b00001000010111100101111000100101;
12'b011011110100: dataB <= 32'b01101001010110011100001100001100;
12'b011011110101: dataB <= 32'b00001111001011111100110110000110;
12'b011011110110: dataB <= 32'b10011001001101111111001010111101;
12'b011011110111: dataB <= 32'b00001000000001011110111110100000;
12'b011011111000: dataB <= 32'b10101110100010011101011100010011;
12'b011011111001: dataB <= 32'b00001110001101110011100100101110;
12'b011011111010: dataB <= 32'b11111001000011000011011111001110;
12'b011011111011: dataB <= 32'b00000011001110100000100011110010;
12'b011011111100: dataB <= 32'b00100011110001100011001010100011;
12'b011011111101: dataB <= 32'b00001001100111011101001010001101;
12'b011011111110: dataB <= 32'b11111010101000001100011001000001;
12'b011011111111: dataB <= 32'b00000100110011011011000010111011;
12'b011100000000: dataB <= 32'b00110010011001100110001100001010;
12'b011100000001: dataB <= 32'b00000111110100101100110001101101;
12'b011100000010: dataB <= 32'b10011100110101111000011000100101;
12'b011100000011: dataB <= 32'b00000001001001010000100000010101;
12'b011100000100: dataB <= 32'b11101011110110101101011101110001;
12'b011100000101: dataB <= 32'b00001111001101100001111010111101;
12'b011100000110: dataB <= 32'b11111011001110110100011000111011;
12'b011100000111: dataB <= 32'b00000001110010100010010110111100;
12'b011100001000: dataB <= 32'b01011010111001010000100100100110;
12'b011100001001: dataB <= 32'b00000100110111011101001101010100;
12'b011100001010: dataB <= 32'b01011010100001100001010010010001;
12'b011100001011: dataB <= 32'b00001001011101101011100110010000;
12'b011100001100: dataB <= 32'b00000000000010110001111010001011;
12'b011100001101: dataB <= 32'b00000000000000000000000000000000;
12'b011100001110: dataB <= 32'b00101000001101010000011000000001;
12'b011100001111: dataB <= 32'b00000110010100100100100100111111;
12'b011100010000: dataB <= 32'b11111100111100010100100010101110;
12'b011100010001: dataB <= 32'b00001000011110101101101111011010;
12'b011100010010: dataB <= 32'b00001100010010011101111011110100;
12'b011100010011: dataB <= 32'b00000101011110011111011000011010;
12'b011100010100: dataB <= 32'b01100000100001000010000110101010;
12'b011100010101: dataB <= 32'b00001011010001110100110100100110;
12'b011100010110: dataB <= 32'b00111010100001111101111001010011;
12'b011100010111: dataB <= 32'b00000111000110100100000110000111;
12'b011100011000: dataB <= 32'b01011100111000101110100100110100;
12'b011100011001: dataB <= 32'b00000111010111110100010101010100;
12'b011100011010: dataB <= 32'b11100110111110110101011110010100;
12'b011100011011: dataB <= 32'b00001011101001100011101010000100;
12'b011100011100: dataB <= 32'b01000111000111001101011111010000;
12'b011100011101: dataB <= 32'b00000111011110101101000000010010;
12'b011100011110: dataB <= 32'b01010001001100110100110101110001;
12'b011100011111: dataB <= 32'b00001011000010011011011001010001;
12'b011100100000: dataB <= 32'b00110101100010100111101111001111;
12'b011100100001: dataB <= 32'b00001000011000011111111010101111;
12'b011100100010: dataB <= 32'b01100100010110011101111101011010;
12'b011100100011: dataB <= 32'b00001000110110110010110101111000;
12'b011100100100: dataB <= 32'b11011010101010000011110111010101;
12'b011100100101: dataB <= 32'b00000110011110110010011001010011;
12'b011100100110: dataB <= 32'b11111000011100001101000001111000;
12'b011100100111: dataB <= 32'b00001000010100011111100110010101;
12'b011100101000: dataB <= 32'b11011010010110100010110111110111;
12'b011100101001: dataB <= 32'b00001110101001111100111100111000;
12'b011100101010: dataB <= 32'b10010010110101010101111011100101;
12'b011100101011: dataB <= 32'b00000011011011011110111001011001;
12'b011100101100: dataB <= 32'b00001010010100010101110011010010;
12'b011100101101: dataB <= 32'b00000010010110010010111100001100;
12'b011100101110: dataB <= 32'b01011110000101010000010101110100;
12'b011100101111: dataB <= 32'b00001000111011101011011100101011;
12'b011100110000: dataB <= 32'b10010010111101110011000110010001;
12'b011100110001: dataB <= 32'b00000110000101011100101100110010;
12'b011100110010: dataB <= 32'b00101101100101011111101100001011;
12'b011100110011: dataB <= 32'b00000011000100010010101110111101;
12'b011100110100: dataB <= 32'b00110000101101010111101000110000;
12'b011100110101: dataB <= 32'b00000001010111011000011110011101;
12'b011100110110: dataB <= 32'b01100100100010111101001110101010;
12'b011100110111: dataB <= 32'b00000011101100010110100110000011;
12'b011100111000: dataB <= 32'b10010011001000011110000101010100;
12'b011100111001: dataB <= 32'b00000101010110100010110000011100;
12'b011100111010: dataB <= 32'b10010101001001110001000011010111;
12'b011100111011: dataB <= 32'b00001001011011111011001001110001;
12'b011100111100: dataB <= 32'b00110001101101110111101001111000;
12'b011100111101: dataB <= 32'b00000100010111100110011010101100;
12'b011100111110: dataB <= 32'b10011000111010010010101011100101;
12'b011100111111: dataB <= 32'b00001010101101110100101000110011;
12'b011101000000: dataB <= 32'b01010010110111010011111011011101;
12'b011101000001: dataB <= 32'b00000011010001011010010100110100;
12'b011101000010: dataB <= 32'b11010010011001001101100110010010;
12'b011101000011: dataB <= 32'b00001000111001101110111000001010;
12'b011101000100: dataB <= 32'b00110011010111010010111111001100;
12'b011101000101: dataB <= 32'b00000001010001011010101011011100;
12'b011101000110: dataB <= 32'b01011101100110011111101100110010;
12'b011101000111: dataB <= 32'b00000110010000011110110010111001;
12'b011101001000: dataB <= 32'b10011000101001111110011101001001;
12'b011101001001: dataB <= 32'b00001001010110101011110100101101;
12'b011101001010: dataB <= 32'b01101011010010011011111011101010;
12'b011101001011: dataB <= 32'b00001110001000111100101010001110;
12'b011101001100: dataB <= 32'b10011001001110010111001100011100;
12'b011101001101: dataB <= 32'b00000110100001011110111110001000;
12'b011101001110: dataB <= 32'b00101010011110100101001100110001;
12'b011101001111: dataB <= 32'b00001101101010110101011101000111;
12'b011101010000: dataB <= 32'b00111000110110111011001110101011;
12'b011101010001: dataB <= 32'b00000011010000011110100011100010;
12'b011101010010: dataB <= 32'b00100111110001100011001001000010;
12'b011101010011: dataB <= 32'b00001000100110011101001010010101;
12'b011101010100: dataB <= 32'b10111000011100001101000111100001;
12'b011101010101: dataB <= 32'b00000101010100011011000010111011;
12'b011101010110: dataB <= 32'b00101110010101110110011011001001;
12'b011101010111: dataB <= 32'b00001000010100101010101101110101;
12'b011101011000: dataB <= 32'b00011010110101100000010111000101;
12'b011101011001: dataB <= 32'b00000000101100001100100100011110;
12'b011101011010: dataB <= 32'b10110001110010110101001101101111;
12'b011101011011: dataB <= 32'b00001110101010100111111011001101;
12'b011101011100: dataB <= 32'b10111101000010110100001010011011;
12'b011101011101: dataB <= 32'b00000010010101011110010110111100;
12'b011101011110: dataB <= 32'b10011010111000111000110011101000;
12'b011101011111: dataB <= 32'b00000101111000011101001101010100;
12'b011101100000: dataB <= 32'b01010110100101010001100010010100;
12'b011101100001: dataB <= 32'b00001010011100101101100010000000;
12'b011101100010: dataB <= 32'b00000000000010101001101001101011;
12'b011101100011: dataB <= 32'b00000000000000000000000000000000;
12'b011101100100: dataB <= 32'b01100010001001000000110110100001;
12'b011101100101: dataB <= 32'b00000110110101100010100101001111;
12'b011101100110: dataB <= 32'b01111100110000010101010010110000;
12'b011101100111: dataB <= 32'b00001001111110110001100111010010;
12'b011101101000: dataB <= 32'b10001000011010101101101100010010;
12'b011101101001: dataB <= 32'b00000110111110100011011000001010;
12'b011101101010: dataB <= 32'b11011110100000111010100110001011;
12'b011101101011: dataB <= 32'b00001011001111110010101100110110;
12'b011101101100: dataB <= 32'b00110110011010000101111001110011;
12'b011101101101: dataB <= 32'b00000110000111011110000110010111;
12'b011101101110: dataB <= 32'b10011100111001000111000101010101;
12'b011101101111: dataB <= 32'b00000111110111101110001101011100;
12'b011101110000: dataB <= 32'b11100110111010111101001110110001;
12'b011101110001: dataB <= 32'b00001011001000100111101010001100;
12'b011101110010: dataB <= 32'b00001001001111010100111111001110;
12'b011101110011: dataB <= 32'b00001000111110101100111000001011;
12'b011101110100: dataB <= 32'b10010011010100110101010110010001;
12'b011101110101: dataB <= 32'b00001001100001011101011001000001;
12'b011101110110: dataB <= 32'b10110111011010111111011111001101;
12'b011101110111: dataB <= 32'b00001000110111100101111011000110;
12'b011101111000: dataB <= 32'b01100000010110101101101110011000;
12'b011101111001: dataB <= 32'b00001001010101110000101101100000;
12'b011101111010: dataB <= 32'b00011000101110000011110111110110;
12'b011101111011: dataB <= 32'b00000111111110101110010001010100;
12'b011101111100: dataB <= 32'b10110100010100010101110010111011;
12'b011101111101: dataB <= 32'b00001000110100100011100110100101;
12'b011101111110: dataB <= 32'b01010110011010011010101000010111;
12'b011101111111: dataB <= 32'b00001101100110111100110100100001;
12'b011110000000: dataB <= 32'b11010010111001100110001010000011;
12'b011110000001: dataB <= 32'b00000100011101011110111001010001;
12'b011110000010: dataB <= 32'b11000110011100100110010011110100;
12'b011110000011: dataB <= 32'b00000011011000010011000100001100;
12'b011110000100: dataB <= 32'b11011000000101000000110110010101;
12'b011110000101: dataB <= 32'b00001010011010101101011000101011;
12'b011110000110: dataB <= 32'b00010011000101101011010110110010;
12'b011110000111: dataB <= 32'b00000101000110011100110000101011;
12'b011110001000: dataB <= 32'b10110001011101110111101011101001;
12'b011110001001: dataB <= 32'b00000010000110010000110011000100;
12'b011110001010: dataB <= 32'b11101110100101101111101000110000;
12'b011110001011: dataB <= 32'b00000010011001010110100010100100;
12'b011110001100: dataB <= 32'b01100010100011000100101101101000;
12'b011110001101: dataB <= 32'b00000011101110010100101001111011;
12'b011110001110: dataB <= 32'b00010011001100101110110101110101;
12'b011110001111: dataB <= 32'b00000101110111100010110000100101;
12'b011110010000: dataB <= 32'b10010111001101011001010100011001;
12'b011110010001: dataB <= 32'b00001010111010111010111101100001;
12'b011110010010: dataB <= 32'b11110101100110001111101010010111;
12'b011110010011: dataB <= 32'b00000101011000100010011010101011;
12'b011110010100: dataB <= 32'b00010110111110001010101010100100;
12'b011110010101: dataB <= 32'b00001010001100110000100000110100;
12'b011110010110: dataB <= 32'b11010010111011010011011100111011;
12'b011110010111: dataB <= 32'b00000011110011010110011000110100;
12'b011110011000: dataB <= 32'b10001110100001010101110110010011;
12'b011110011001: dataB <= 32'b00001001111000101110110000001011;
12'b011110011010: dataB <= 32'b10110101001111001010011110101001;
12'b011110011011: dataB <= 32'b00000001110100011000101111011011;
12'b011110011100: dataB <= 32'b00100001100110110111011101010000;
12'b011110011101: dataB <= 32'b00000110010001011100110010101001;
12'b011110011110: dataB <= 32'b00010110101110001110011100000111;
12'b011110011111: dataB <= 32'b00001001110110110001110000111110;
12'b011110100000: dataB <= 32'b00101101001010011011101011001001;
12'b011110100001: dataB <= 32'b00001101100110111000100010011110;
12'b011110100010: dataB <= 32'b10011011010010100110111101011010;
12'b011110100011: dataB <= 32'b00000101000001011110111101110000;
12'b011110100100: dataB <= 32'b10100110011010101100111100101111;
12'b011110100101: dataB <= 32'b00001101001000111001010001010111;
12'b011110100110: dataB <= 32'b10110110101110110010101110001001;
12'b011110100111: dataB <= 32'b00000011010010011010100111011001;
12'b011110101000: dataB <= 32'b00101011101101011011010111100010;
12'b011110101001: dataB <= 32'b00000111100110011111001010010101;
12'b011110101010: dataB <= 32'b00110100010100010101110110000001;
12'b011110101011: dataB <= 32'b00000101110101011011000110111011;
12'b011110101100: dataB <= 32'b01101000001110000110011010101000;
12'b011110101101: dataB <= 32'b00001000110100101000101001111101;
12'b011110101110: dataB <= 32'b11011010111001010000100110000101;
12'b011110101111: dataB <= 32'b00000000101111001010101100101110;
12'b011110110000: dataB <= 32'b00110101101010111100111101101101;
12'b011110110001: dataB <= 32'b00001110000111101101110111010101;
12'b011110110010: dataB <= 32'b00111100111010110011101011011010;
12'b011110110011: dataB <= 32'b00000010110111011010010111000100;
12'b011110110100: dataB <= 32'b11011010111100101001010011001001;
12'b011110110101: dataB <= 32'b00000110111001011111010001011100;
12'b011110110110: dataB <= 32'b01010100101001001001110010110110;
12'b011110110111: dataB <= 32'b00001011011011110001011001101000;
12'b011110111000: dataB <= 32'b00000000000010011001011001001010;
12'b011110111001: dataB <= 32'b00000000000000000000000000000000;
12'b011110111010: dataB <= 32'b10011110001000101001010101100001;
12'b011110111011: dataB <= 32'b00000111010101011110100001100111;
12'b011110111100: dataB <= 32'b11111010100100100101110010110011;
12'b011110111101: dataB <= 32'b00001011011101110101100011000001;
12'b011110111110: dataB <= 32'b01000100100110110101011100010000;
12'b011110111111: dataB <= 32'b00001000011110100101011000001011;
12'b011111000000: dataB <= 32'b01011010100000110011000101101100;
12'b011111000001: dataB <= 32'b00001011001110110000100101001111;
12'b011111000010: dataB <= 32'b11110010010010010101111001110010;
12'b011111000011: dataB <= 32'b00000101001000011000000110100110;
12'b011111000100: dataB <= 32'b11011100111001010111100101110110;
12'b011111000101: dataB <= 32'b00001000110111101010000101011100;
12'b011111000110: dataB <= 32'b11100110111010111100101110101111;
12'b011111000111: dataB <= 32'b00001010000111101011100110001100;
12'b011111001000: dataB <= 32'b11001011010111010100011110101011;
12'b011111001001: dataB <= 32'b00001010011110101100110100001011;
12'b011111001010: dataB <= 32'b00010101011001000101110110010010;
12'b011111001011: dataB <= 32'b00001000000001100001011100110010;
12'b011111001100: dataB <= 32'b01111001010011001110111110101010;
12'b011111001101: dataB <= 32'b00001001110111101001111011010110;
12'b011111001110: dataB <= 32'b10011010010110110101011110110110;
12'b011111001111: dataB <= 32'b00001001110101101110100101001000;
12'b011111010000: dataB <= 32'b01010110110010000011111000010110;
12'b011111010001: dataB <= 32'b00001001011110101010001101010100;
12'b011111010010: dataB <= 32'b01110000001100100110010100011100;
12'b011111010011: dataB <= 32'b00001001010100100111100110101101;
12'b011111010100: dataB <= 32'b00010010011110010010101001010111;
12'b011111010101: dataB <= 32'b00001101000100111010101000011010;
12'b011111010110: dataB <= 32'b01010001000001110110001001000011;
12'b011111010111: dataB <= 32'b00000101111110011110111001000010;
12'b011111011000: dataB <= 32'b10000100100100110110110100010110;
12'b011111011001: dataB <= 32'b00000011111010010011001000010101;
12'b011111011010: dataB <= 32'b10010010001000101001010110110101;
12'b011111011011: dataB <= 32'b00001011011001101111010000101100;
12'b011111011100: dataB <= 32'b10010011001001101011010110110010;
12'b011111011101: dataB <= 32'b00000100000111011010110000101011;
12'b011111011110: dataB <= 32'b00110011010110001111101010101000;
12'b011111011111: dataB <= 32'b00000001001001010000111011000100;
12'b011111100000: dataB <= 32'b10101010100010000111101000110000;
12'b011111100001: dataB <= 32'b00000011011011010010100110100100;
12'b011111100010: dataB <= 32'b01011110011111000100001101000101;
12'b011111100011: dataB <= 32'b00000011010000010010101101111011;
12'b011111100100: dataB <= 32'b10010101010001000111000110010110;
12'b011111100101: dataB <= 32'b00000110110111100000110000101101;
12'b011111100110: dataB <= 32'b11011001010001001001100100111010;
12'b011111100111: dataB <= 32'b00001011111001111010110101010001;
12'b011111101000: dataB <= 32'b10111001011110100111101011010110;
12'b011111101001: dataB <= 32'b00000110011001011110010110101011;
12'b011111101010: dataB <= 32'b10010111000010000010101001100011;
12'b011111101011: dataB <= 32'b00001001101011101100011000110100;
12'b011111101100: dataB <= 32'b01010001000011001010111101111001;
12'b011111101101: dataB <= 32'b00000100010101010010011100111101;
12'b011111101110: dataB <= 32'b01001100101001100110000110110011;
12'b011111101111: dataB <= 32'b00001010110111101100101100001100;
12'b011111110000: dataB <= 32'b00110101000110111001111110000111;
12'b011111110001: dataB <= 32'b00000010010110010110110011010011;
12'b011111110010: dataB <= 32'b11100101100111000110111101001110;
12'b011111110011: dataB <= 32'b00000110010001011100110010011000;
12'b011111110100: dataB <= 32'b10010100110010011110011011100101;
12'b011111110101: dataB <= 32'b00001010010101110101101001000110;
12'b011111110110: dataB <= 32'b11101101000110011011101010001000;
12'b011111110111: dataB <= 32'b00001100100100110100010110101101;
12'b011111111000: dataB <= 32'b10011101010010110110101110011000;
12'b011111111001: dataB <= 32'b00000100000011011110111101100000;
12'b011111111010: dataB <= 32'b10100010011010101100101100101101;
12'b011111111011: dataB <= 32'b00001100000110111001001001101111;
12'b011111111100: dataB <= 32'b00110100100110101010011101000111;
12'b011111111101: dataB <= 32'b00000011110100011000100111001001;
12'b011111111110: dataB <= 32'b11110001100101011011100110100010;
12'b011111111111: dataB <= 32'b00000110100110011111001010011100;
12'b100000000000: dataB <= 32'b11110000001100100110010100100010;
12'b100000000001: dataB <= 32'b00000110010110011011000110110010;
12'b100000000010: dataB <= 32'b01100100001110010110011001100111;
12'b100000000011: dataB <= 32'b00001001010100100110100110000101;
12'b100000000100: dataB <= 32'b00011010111000111000110101000110;
12'b100000000101: dataB <= 32'b00000000110010001010110101000111;
12'b100000000110: dataB <= 32'b10111001100010111100011101001011;
12'b100000000111: dataB <= 32'b00001101000101110001110011010100;
12'b100000001000: dataB <= 32'b10111010101110110011011100011000;
12'b100000001001: dataB <= 32'b00000011111001010110011011000011;
12'b100000001010: dataB <= 32'b00011010111100011001110010101011;
12'b100000001011: dataB <= 32'b00000111111001100001010001100101;
12'b100000001100: dataB <= 32'b10010010101100111010010011111000;
12'b100000001101: dataB <= 32'b00001100111001110011010001010000;
12'b100000001110: dataB <= 32'b00000000000010001001011000101010;
12'b100000001111: dataB <= 32'b00000000000000000000000000000000;
12'b100000010000: dataB <= 32'b11000101000000101110100000110100;
12'b100000010001: dataB <= 32'b00001010110001010001000011110100;
12'b100000010010: dataB <= 32'b11010010001010111110111001111010;
12'b100000010011: dataB <= 32'b00001110101001110000010100111001;
12'b100000010100: dataB <= 32'b10010011110110101010011000000111;
12'b100000010101: dataB <= 32'b00001111001111101100110101101111;
12'b100000010110: dataB <= 32'b10010001001001100110010110010100;
12'b100000010111: dataB <= 32'b00000111001001010010011111101101;
12'b100000011000: dataB <= 32'b11001000011010111011011001001100;
12'b100000011001: dataB <= 32'b00000100010101000011001111011010;
12'b100000011010: dataB <= 32'b00011101000111110101011011010100;
12'b100000011011: dataB <= 32'b00001011101110000010101010011101;
12'b100000011100: dataB <= 32'b10011100110010010010000111100010;
12'b100000011101: dataB <= 32'b00000011101011110010101010011011;
12'b100000011110: dataB <= 32'b10101011101010001001010101100010;
12'b100000011111: dataB <= 32'b00001111001011011010100101111111;
12'b100000100000: dataB <= 32'b01101101010110111101111001010011;
12'b100000100001: dataB <= 32'b00000000101111101110111101000110;
12'b100000100010: dataB <= 32'b01101000001111011001100101000010;
12'b100000100011: dataB <= 32'b00001011101100111100101111001001;
12'b100000100100: dataB <= 32'b10001011001010101010011011000010;
12'b100000100101: dataB <= 32'b00001010101100010010100000010101;
12'b100000100110: dataB <= 32'b01011001010001111011111011001111;
12'b100000100111: dataB <= 32'b00001111001101000110101010001101;
12'b100000101000: dataB <= 32'b10000110011111001110111110010111;
12'b100000101001: dataB <= 32'b00001010001101110010110010101010;
12'b100000101010: dataB <= 32'b00001111011001010011011011101101;
12'b100000101011: dataB <= 32'b00000010000101010100001001000111;
12'b100000101100: dataB <= 32'b11100001011111000100010001101101;
12'b100000101101: dataB <= 32'b00001111010100011101000001001101;
12'b100000101110: dataB <= 32'b01010011110111011110011011010111;
12'b100000101111: dataB <= 32'b00001101011000100101011010110111;
12'b100000110000: dataB <= 32'b10000101011000101110101010110010;
12'b100000110001: dataB <= 32'b00001100101001101000100010010110;
12'b100000110010: dataB <= 32'b10100101011001101100101001010010;
12'b100000110011: dataB <= 32'b00000011110111011001001001110110;
12'b100000110100: dataB <= 32'b11101010011011110011100100001010;
12'b100000110101: dataB <= 32'b00000100111101011101011110000001;
12'b100000110110: dataB <= 32'b11010000101011110011111000001110;
12'b100000110111: dataB <= 32'b00001101111001010011011010010010;
12'b100000111000: dataB <= 32'b00001111000010000001110010100101;
12'b100000111001: dataB <= 32'b00001000011001010111011001101100;
12'b100000111010: dataB <= 32'b10101001010111100101111011010011;
12'b100000111011: dataB <= 32'b00001011110010011000111110110110;
12'b100000111100: dataB <= 32'b01101001001100110101101101010110;
12'b100000111101: dataB <= 32'b00001100101000011010001000111101;
12'b100000111110: dataB <= 32'b10101110001111110010111011001001;
12'b100000111111: dataB <= 32'b00001100110011001011000001110010;
12'b100001000000: dataB <= 32'b01100001010001010011110001101100;
12'b100001000001: dataB <= 32'b00000101101100001100100110010110;
12'b100001000010: dataB <= 32'b00100001011101011001101100100100;
12'b100001000011: dataB <= 32'b00001010110111001111011010101110;
12'b100001000100: dataB <= 32'b10010101100111000100111001110010;
12'b100001000101: dataB <= 32'b00001011101010010110100110001111;
12'b100001000110: dataB <= 32'b01100010010100111010000011100011;
12'b100001000111: dataB <= 32'b00001011011011011001010001100001;
12'b100001001000: dataB <= 32'b00110010110111011001110111000101;
12'b100001001001: dataB <= 32'b00001000110011011001000100011011;
12'b100001001010: dataB <= 32'b11011001010111001011000010101000;
12'b100001001011: dataB <= 32'b00001010101011110100010111010101;
12'b100001001100: dataB <= 32'b10100010100101110011000100001011;
12'b100001001101: dataB <= 32'b00000010000110001010010110111010;
12'b100001001110: dataB <= 32'b11101001000111010010011100000011;
12'b100001001111: dataB <= 32'b00000001110111011111000000010100;
12'b100001010000: dataB <= 32'b10001100111010010010100110100110;
12'b100001010001: dataB <= 32'b00000011000111100100001111110100;
12'b100001010010: dataB <= 32'b10010010010101001010100011100101;
12'b100001010011: dataB <= 32'b00001010011000010011001100100001;
12'b100001010100: dataB <= 32'b00110010011101110101000001010010;
12'b100001010101: dataB <= 32'b00000011010010100101000010011011;
12'b100001010110: dataB <= 32'b01000110011111001110110001010110;
12'b100001010111: dataB <= 32'b00001011010011100011001001011010;
12'b100001011000: dataB <= 32'b11000110110111001011010011101100;
12'b100001011001: dataB <= 32'b00001010001101010010110010101011;
12'b100001011010: dataB <= 32'b11011101001000011110000011010101;
12'b100001011011: dataB <= 32'b00001001011110011011101011100101;
12'b100001011100: dataB <= 32'b01110000001110001010000101100101;
12'b100001011101: dataB <= 32'b00000010100101111000011110010001;
12'b100001011110: dataB <= 32'b11010110001001101010011100000111;
12'b100001011111: dataB <= 32'b00001100111000001101010001110001;
12'b100001100000: dataB <= 32'b11011111001000111111000101111010;
12'b100001100001: dataB <= 32'b00001100110000101000111110100100;
12'b100001100010: dataB <= 32'b01010111011001001110001100011000;
12'b100001100011: dataB <= 32'b00001100100110101000011000010101;
12'b100001100100: dataB <= 32'b00000000000000101011100101001110;
12'b100001100101: dataB <= 32'b00000000000000000000000000000000;
12'b100001100110: dataB <= 32'b10000100111000011101110000110010;
12'b100001100111: dataB <= 32'b00001010110010010010111011101101;
12'b100001101000: dataB <= 32'b01011000000110101111011000011010;
12'b100001101001: dataB <= 32'b00001111001100110010011101001001;
12'b100001101010: dataB <= 32'b10001101101110110010101001000111;
12'b100001101011: dataB <= 32'b00001111010010101100111001010111;
12'b100001101100: dataB <= 32'b01010001000001010110000101110011;
12'b100001101101: dataB <= 32'b00000111101001010110011011011110;
12'b100001101110: dataB <= 32'b01001100010010111011111001101100;
12'b100001101111: dataB <= 32'b00000011110011000011000011100011;
12'b100001110000: dataB <= 32'b00011101000111100101111010110101;
12'b100001110001: dataB <= 32'b00001011110000000110100010010101;
12'b100001110010: dataB <= 32'b10011100110010100010001000100010;
12'b100001110011: dataB <= 32'b00000100001001110100110010011011;
12'b100001110100: dataB <= 32'b10100111101110011001010111000001;
12'b100001110101: dataB <= 32'b00001111001110011100100101100111;
12'b100001110110: dataB <= 32'b11101011011010101110011000110011;
12'b100001110111: dataB <= 32'b00000000101100101101000100110101;
12'b100001111000: dataB <= 32'b11101100010011101010000110100001;
12'b100001111001: dataB <= 32'b00001011101110111100110111010001;
12'b100001111010: dataB <= 32'b11001010111110110010101100000011;
12'b100001111011: dataB <= 32'b00001010101101010110011100001100;
12'b100001111100: dataB <= 32'b01010111001101111011111011010000;
12'b100001111101: dataB <= 32'b00001111010000001000100010000101;
12'b100001111110: dataB <= 32'b11001010010110111111011101111010;
12'b100001111111: dataB <= 32'b00001010001110110010111010110010;
12'b100010000000: dataB <= 32'b11001101010001010011001011101111;
12'b100010000001: dataB <= 32'b00000011000100011010000100101110;
12'b100010000010: dataB <= 32'b01011101011011000100110001101011;
12'b100010000011: dataB <= 32'b00001110110111011101000000111101;
12'b100010000100: dataB <= 32'b10001111110011001110111010011000;
12'b100010000101: dataB <= 32'b00001100011001100011011010011111;
12'b100010000110: dataB <= 32'b10000011001100011101111010110011;
12'b100010000111: dataB <= 32'b00001101001011101100100101111110;
12'b100010001000: dataB <= 32'b10100011011001101100101001010010;
12'b100010001001: dataB <= 32'b00000011010101011001000101100110;
12'b100010001010: dataB <= 32'b11101110011111110100010100101000;
12'b100010001011: dataB <= 32'b00000011011011011001011110010001;
12'b100010001100: dataB <= 32'b11010010100011110100101000001110;
12'b100010001101: dataB <= 32'b00001100111011010001010010011010;
12'b100010001110: dataB <= 32'b00010000111010010001110100000100;
12'b100010001111: dataB <= 32'b00000111011000010101010101101100;
12'b100010010000: dataB <= 32'b11100111011011011110101010110100;
12'b100010010001: dataB <= 32'b00001011110100011000111010100110;
12'b100010010010: dataB <= 32'b11100111010000101101001100110111;
12'b100010010011: dataB <= 32'b00001101001010011110001000110100;
12'b100010010100: dataB <= 32'b10110010010111110011101011101011;
12'b100010010101: dataB <= 32'b00001100010101001100111001111010;
12'b100010010110: dataB <= 32'b01011111010001010011100010001010;
12'b100010010111: dataB <= 32'b00000110001011010000011110000110;
12'b100010011000: dataB <= 32'b01011101011001101001011101100110;
12'b100010011001: dataB <= 32'b00001001111000001101010010011110;
12'b100010011010: dataB <= 32'b10010001100010111101011001110011;
12'b100010011011: dataB <= 32'b00001100001100011000100001110111;
12'b100010011100: dataB <= 32'b00100110010101001001100100100010;
12'b100010011101: dataB <= 32'b00001010011100010111001101110001;
12'b100010011110: dataB <= 32'b10110010111111101010011000000101;
12'b100010011111: dataB <= 32'b00001000110011011001000100100010;
12'b100010100000: dataB <= 32'b00010111010011001011100011100111;
12'b100010100001: dataB <= 32'b00001011001100111000011111000110;
12'b100010100010: dataB <= 32'b00100100100101110011000100101001;
12'b100010100011: dataB <= 32'b00000011000100010000001111000011;
12'b100010100100: dataB <= 32'b01101001001011011010111101000101;
12'b100010100101: dataB <= 32'b00000000110101011111000000010100;
12'b100010100110: dataB <= 32'b01001100110010011010100111100110;
12'b100010100111: dataB <= 32'b00000100000101101000001111110101;
12'b100010101000: dataB <= 32'b00010110010001010010010100100011;
12'b100010101001: dataB <= 32'b00001001011001010011001000110001;
12'b100010101010: dataB <= 32'b01110110101001101101000001010000;
12'b100010101011: dataB <= 32'b00000011010000100101000010100011;
12'b100010101100: dataB <= 32'b00001010010110111111010000110011;
12'b100010101101: dataB <= 32'b00001010110100100011001001100010;
12'b100010101110: dataB <= 32'b00000110101111001011110100001010;
12'b100010101111: dataB <= 32'b00001010001110010100101110101100;
12'b100010110000: dataB <= 32'b10011101001000010101010010110011;
12'b100010110001: dataB <= 32'b00000111111110010111101011011110;
12'b100010110010: dataB <= 32'b01110100010110011010000110100100;
12'b100010110011: dataB <= 32'b00000011100011111010100110100001;
12'b100010110100: dataB <= 32'b11011100000101110010011101001001;
12'b100010110101: dataB <= 32'b00001011111010001011001010000001;
12'b100010110110: dataB <= 32'b00011111001000101110100100111001;
12'b100010110111: dataB <= 32'b00001100110010101001000010011101;
12'b100010111000: dataB <= 32'b10010101010100111101101011011010;
12'b100010111001: dataB <= 32'b00001101101001101100011100001100;
12'b100010111010: dataB <= 32'b00000000000000101011000101001101;
12'b100010111011: dataB <= 32'b00000000000000000000000000000000;
12'b100010111100: dataB <= 32'b00000110101100001101010000101111;
12'b100010111101: dataB <= 32'b00001010010011010010110111100110;
12'b100010111110: dataB <= 32'b00011110000110010111010111011010;
12'b100010111111: dataB <= 32'b00001111001111110110100101011001;
12'b100011000000: dataB <= 32'b00001001100110111011001010001000;
12'b100011000001: dataB <= 32'b00001111010101101101000001000111;
12'b100011000010: dataB <= 32'b11010000111101000101110101010010;
12'b100011000011: dataB <= 32'b00001000101001011010010111001110;
12'b100011000100: dataB <= 32'b11010000001010111100001001101101;
12'b100011000101: dataB <= 32'b00000011010001000010110111100011;
12'b100011000110: dataB <= 32'b01011101000111010110101010010110;
12'b100011000111: dataB <= 32'b00001011110001001010010110001101;
12'b100011001000: dataB <= 32'b11011110110010101010011010000011;
12'b100011001001: dataB <= 32'b00000100101000110100111010011011;
12'b100011001010: dataB <= 32'b01100011110010101001101000000001;
12'b100011001011: dataB <= 32'b00001111010001100000100101001111;
12'b100011001100: dataB <= 32'b01100111011110011110011000110100;
12'b100011001101: dataB <= 32'b00000001001001101101001000101101;
12'b100011001110: dataB <= 32'b10110000010111110010110111100001;
12'b100011001111: dataB <= 32'b00001100001111111101000011100010;
12'b100011010000: dataB <= 32'b00001010110110111011001101000101;
12'b100011010001: dataB <= 32'b00001011001110011010011000001100;
12'b100011010010: dataB <= 32'b01010101001001111011111010110001;
12'b100011010011: dataB <= 32'b00001111010011001100011001111101;
12'b100011010100: dataB <= 32'b01001110001110100111101100011100;
12'b100011010101: dataB <= 32'b00001010001111110011000010111011;
12'b100011010110: dataB <= 32'b00001011001001011010111011110000;
12'b100011010111: dataB <= 32'b00000100100010011110000100011110;
12'b100011011000: dataB <= 32'b00011011011010111101010010101000;
12'b100011011001: dataB <= 32'b00001101111001011101000000110101;
12'b100011011010: dataB <= 32'b10001011101010111111011001011001;
12'b100011011011: dataB <= 32'b00001011011011011111011010000111;
12'b100011011100: dataB <= 32'b10000011000000001101011010010100;
12'b100011011101: dataB <= 32'b00001101101110101110101001101110;
12'b100011011110: dataB <= 32'b01011111011001100100011000110011;
12'b100011011111: dataB <= 32'b00000010110011010111000101010110;
12'b100011100000: dataB <= 32'b00110010100111110101000101100111;
12'b100011100001: dataB <= 32'b00000010011001010111011010100010;
12'b100011100010: dataB <= 32'b00010110011111110101011000001110;
12'b100011100011: dataB <= 32'b00001011111101001111001110100011;
12'b100011100100: dataB <= 32'b11010000110110100010000101000010;
12'b100011100101: dataB <= 32'b00000110011000010011010001101011;
12'b100011100110: dataB <= 32'b00100101011011000111001010010101;
12'b100011100111: dataB <= 32'b00001011010101011000111010010111;
12'b100011101000: dataB <= 32'b01100101010100100100011011111001;
12'b100011101001: dataB <= 32'b00001101101101100100001000110100;
12'b100011101010: dataB <= 32'b10110110011111110100011100001100;
12'b100011101011: dataB <= 32'b00001011110111001100110010000010;
12'b100011101100: dataB <= 32'b01011101001101010011010010101000;
12'b100011101101: dataB <= 32'b00000110101010010100010101110110;
12'b100011101110: dataB <= 32'b01011011011001111001011110101001;
12'b100011101111: dataB <= 32'b00001000111001001011001010001110;
12'b100011110000: dataB <= 32'b10001101011010110101101001010011;
12'b100011110001: dataB <= 32'b00001100101110011100100001011111;
12'b100011110010: dataB <= 32'b00101010011001011001010110000001;
12'b100011110011: dataB <= 32'b00001000111101010101001010000001;
12'b100011110100: dataB <= 32'b00110011000111110011001001000110;
12'b100011110101: dataB <= 32'b00001000010011011001000000101010;
12'b100011110110: dataB <= 32'b10010101001111001100000100100101;
12'b100011110111: dataB <= 32'b00001011001101111010101010110110;
12'b100011111000: dataB <= 32'b10101000101001111011000101001000;
12'b100011111001: dataB <= 32'b00000100000011010100000111001011;
12'b100011111010: dataB <= 32'b10100111001111100011011110000111;
12'b100011111011: dataB <= 32'b00000000110010011111000000010011;
12'b100011111100: dataB <= 32'b11001110101010100010111000100110;
12'b100011111101: dataB <= 32'b00000101000100101110010111100101;
12'b100011111110: dataB <= 32'b11011010001101100010000101100010;
12'b100011111111: dataB <= 32'b00001000011001010001000001000000;
12'b100100000000: dataB <= 32'b01111000110001100100110001001101;
12'b100100000001: dataB <= 32'b00000011001110100101000110100011;
12'b100100000010: dataB <= 32'b00001110001110100111100000110000;
12'b100100000011: dataB <= 32'b00001010010101100001001001110010;
12'b100100000100: dataB <= 32'b01001010100011001100010100101001;
12'b100100000101: dataB <= 32'b00001010001111010110101010100100;
12'b100100000110: dataB <= 32'b00011011001000001100110010110001;
12'b100100000111: dataB <= 32'b00000110011110010011100111000111;
12'b100100001000: dataB <= 32'b10111000011110100010010111100100;
12'b100100001001: dataB <= 32'b00000101000010111100110010110001;
12'b100100001010: dataB <= 32'b00100000000110000010011101101011;
12'b100100001011: dataB <= 32'b00001010111011001011000010010010;
12'b100100001100: dataB <= 32'b01011101001000011110000100011000;
12'b100100001101: dataB <= 32'b00001100010100100111000110010101;
12'b100100001110: dataB <= 32'b11010011010000110101011010011011;
12'b100100001111: dataB <= 32'b00001110001011110000100100001011;
12'b100100010000: dataB <= 32'b00000000000000110010100101101100;
12'b100100010001: dataB <= 32'b00000000000000000000000000000000;
12'b100100010010: dataB <= 32'b10001000100100001100100000101100;
12'b100100010011: dataB <= 32'b00001010010100010010110011010110;
12'b100100010100: dataB <= 32'b00100100000101111111100110011010;
12'b100100010101: dataB <= 32'b00001111010010111000101101110001;
12'b100100010110: dataB <= 32'b10000101011111000011011010101001;
12'b100100010111: dataB <= 32'b00001110010111101101000100101110;
12'b100100011000: dataB <= 32'b01010000110100111101010101010001;
12'b100100011001: dataB <= 32'b00001001001010011110010110111111;
12'b100100011010: dataB <= 32'b10010110000110111100101010001110;
12'b100100011011: dataB <= 32'b00000011010000000010101011100100;
12'b100100011100: dataB <= 32'b01011011000011000111001001010111;
12'b100100011101: dataB <= 32'b00001011010010001110001110000101;
12'b100100011110: dataB <= 32'b00100000110010110010111011000100;
12'b100100011111: dataB <= 32'b00000101100111110101000110011100;
12'b100100100000: dataB <= 32'b00011111110010110001111001100010;
12'b100100100001: dataB <= 32'b00001111010100100010100100111111;
12'b100100100010: dataB <= 32'b11100101100010001110101000010100;
12'b100100100011: dataB <= 32'b00000001100111101101001100100100;
12'b100100100100: dataB <= 32'b00110100011111110011101001000001;
12'b100100100101: dataB <= 32'b00001011110001111101001111101011;
12'b100100100110: dataB <= 32'b01001100101111000011011110001000;
12'b100100100111: dataB <= 32'b00001011010000011110011000001011;
12'b100100101000: dataB <= 32'b01010101000101111011111010110011;
12'b100100101001: dataB <= 32'b00001110110110010000010001110101;
12'b100100101010: dataB <= 32'b10010100001010001111101011011101;
12'b100100101011: dataB <= 32'b00001010010000110011001010111011;
12'b100100101100: dataB <= 32'b10001011000001100010101011110010;
12'b100100101101: dataB <= 32'b00000110000001100100000100010101;
12'b100100101110: dataB <= 32'b10011001011010110101100011000110;
12'b100100101111: dataB <= 32'b00001100111011011101000000110100;
12'b100100110000: dataB <= 32'b10000111011110100111101000011001;
12'b100100110001: dataB <= 32'b00001010011100011101011001101111;
12'b100100110010: dataB <= 32'b01000010110100001100101001110101;
12'b100100110011: dataB <= 32'b00001101110000110000110001011110;
12'b100100110100: dataB <= 32'b00011101011001100100011000110011;
12'b100100110101: dataB <= 32'b00000010010001010111000001001110;
12'b100100110110: dataB <= 32'b01110100101111101101110110000111;
12'b100100110111: dataB <= 32'b00000001010111010101010110101010;
12'b100100111000: dataB <= 32'b01011000011111100101111000101110;
12'b100100111001: dataB <= 32'b00001010011110001101000110100011;
12'b100100111010: dataB <= 32'b11010010101110101010010110100010;
12'b100100111011: dataB <= 32'b00000101110111010001001001101011;
12'b100100111100: dataB <= 32'b00100001011110110111011001110110;
12'b100100111101: dataB <= 32'b00001010010110011000110101111111;
12'b100100111110: dataB <= 32'b11100011010100100011111010111010;
12'b100100111111: dataB <= 32'b00001110001111101010001100110011;
12'b100101000000: dataB <= 32'b10111000100111110101001100101110;
12'b100101000001: dataB <= 32'b00001010111000001110101010001010;
12'b100101000010: dataB <= 32'b00011101001101011011000011100110;
12'b100101000011: dataB <= 32'b00000111001010011000010101100110;
12'b100101000100: dataB <= 32'b01011001011010001001011111001011;
12'b100101000101: dataB <= 32'b00001000011001001011000001111110;
12'b100101000110: dataB <= 32'b01001011010010101110001000110100;
12'b100101000111: dataB <= 32'b00001100101111011110100001000111;
12'b100101001000: dataB <= 32'b01101100011101101001000111100001;
12'b100101001001: dataB <= 32'b00000111111101010101000110010001;
12'b100101001010: dataB <= 32'b10110001001111110011111010000111;
12'b100101001011: dataB <= 32'b00000111110011011000111100111001;
12'b100101001100: dataB <= 32'b11010011001011001100100101100100;
12'b100101001101: dataB <= 32'b00001011101111111100110110100110;
12'b100101001110: dataB <= 32'b11101010101110000011000110000111;
12'b100101001111: dataB <= 32'b00000101100001011010000111001011;
12'b100101010000: dataB <= 32'b11100111001111100100001110101010;
12'b100101010001: dataB <= 32'b00000000101111011111000000010010;
12'b100101010010: dataB <= 32'b10010000100010101011001001100111;
12'b100101010011: dataB <= 32'b00000110100011110010011011010110;
12'b100101010100: dataB <= 32'b01100000001101101001110111000001;
12'b100101010101: dataB <= 32'b00000111011001010000111101011000;
12'b100101010110: dataB <= 32'b10111000111001100100110001101010;
12'b100101010111: dataB <= 32'b00000011101100100101000110100011;
12'b100101011000: dataB <= 32'b00010100001010001111100000101101;
12'b100101011001: dataB <= 32'b00001001110110100001001001111010;
12'b100101011010: dataB <= 32'b10001100011011000100110101000111;
12'b100101011011: dataB <= 32'b00001010010000011000100110100100;
12'b100101011100: dataB <= 32'b01011011000100001100000010101110;
12'b100101011101: dataB <= 32'b00000100111101010001011110110111;
12'b100101011110: dataB <= 32'b00111010101010101010101000100100;
12'b100101011111: dataB <= 32'b00000110100001111100111110111010;
12'b100101100000: dataB <= 32'b00100110001010001010011101101110;
12'b100101100001: dataB <= 32'b00001001011100001010111010011010;
12'b100101100010: dataB <= 32'b01011101001000010101010011010110;
12'b100101100011: dataB <= 32'b00001011110110100111000110001101;
12'b100101100100: dataB <= 32'b01010001001000101100111000111011;
12'b100101100101: dataB <= 32'b00001110101101110010101000001011;
12'b100101100110: dataB <= 32'b00000000000000111010010101101011;
12'b100101100111: dataB <= 32'b00000000000000000000000000000000;
12'b100101101000: dataB <= 32'b00001100011100001011110001001001;
12'b100101101001: dataB <= 32'b00001001110101010100101110111111;
12'b100101101010: dataB <= 32'b11101000000101101111010101011001;
12'b100101101011: dataB <= 32'b00001111010101111000111010000000;
12'b100101101100: dataB <= 32'b00000011010011000011111011001010;
12'b100101101101: dataB <= 32'b00001101011010101101001000011110;
12'b100101101110: dataB <= 32'b10010010110000110101000101010000;
12'b100101101111: dataB <= 32'b00001001101010100010010110100111;
12'b100101110000: dataB <= 32'b00011100000110110100111010001111;
12'b100101110001: dataB <= 32'b00000011001110000110100011011101;
12'b100101110010: dataB <= 32'b01011011000010110111011000110111;
12'b100101110011: dataB <= 32'b00001010110100010010001001111101;
12'b100101110100: dataB <= 32'b01100010110010111011001100000110;
12'b100101110101: dataB <= 32'b00000110100110110101001110011100;
12'b100101110110: dataB <= 32'b10011001101111000010011011000011;
12'b100101110111: dataB <= 32'b00001110110111100100100100101110;
12'b100101111000: dataB <= 32'b00100001100001111110100111110100;
12'b100101111001: dataB <= 32'b00000010100101101011010000011100;
12'b100101111010: dataB <= 32'b11110110101011110100011010100010;
12'b100101111011: dataB <= 32'b00001011110010111011011011101011;
12'b100101111100: dataB <= 32'b11001110101011000011111111001010;
12'b100101111101: dataB <= 32'b00001011010001100000011000001010;
12'b100101111110: dataB <= 32'b00010101000001111011111010010100;
12'b100101111111: dataB <= 32'b00001110011000010100001101101101;
12'b100110000000: dataB <= 32'b00011010000101110111101001111110;
12'b100110000001: dataB <= 32'b00001010010001110001010010111100;
12'b100110000010: dataB <= 32'b11001010111001101010101011010011;
12'b100110000011: dataB <= 32'b00000111100001101010001000001100;
12'b100110000100: dataB <= 32'b00010111010110100101110100000101;
12'b100110000101: dataB <= 32'b00001011111101011100111100110100;
12'b100110000110: dataB <= 32'b10000011010110001111100111111001;
12'b100110000111: dataB <= 32'b00001000111100011011011001010111;
12'b100110001000: dataB <= 32'b00000010101000001011111001010101;
12'b100110001001: dataB <= 32'b00001101110010110000111001010110;
12'b100110001010: dataB <= 32'b10011011011001100100001000010011;
12'b100110001011: dataB <= 32'b00000010001110010110111100111101;
12'b100110001100: dataB <= 32'b10110100110111011110010111000110;
12'b100110001101: dataB <= 32'b00000000110100010011010010110010;
12'b100110001110: dataB <= 32'b10011100011011010110101000101110;
12'b100110001111: dataB <= 32'b00001000111110001100111110101011;
12'b100110010000: dataB <= 32'b11010100101010110010100111100001;
12'b100110010001: dataB <= 32'b00000100110110010001000101101011;
12'b100110010010: dataB <= 32'b00011111011110011111101001010111;
12'b100110010011: dataB <= 32'b00001001110111011010110001101111;
12'b100110010100: dataB <= 32'b01100001010100100011011001111011;
12'b100110010101: dataB <= 32'b00001101110001101110010000110011;
12'b100110010110: dataB <= 32'b11111010110011101101111100110000;
12'b100110010111: dataB <= 32'b00001010011001010000100010010010;
12'b100110011000: dataB <= 32'b00011011001101100010110100100100;
12'b100110011001: dataB <= 32'b00000111101010011100010001010110;
12'b100110011010: dataB <= 32'b01010111010110011001101111001110;
12'b100110011011: dataB <= 32'b00000111011001001010111001101110;
12'b100110011100: dataB <= 32'b11001011001010011110001000010100;
12'b100110011101: dataB <= 32'b00001100110001100010100000110110;
12'b100110011110: dataB <= 32'b01110000100101111001001001000001;
12'b100110011111: dataB <= 32'b00000110011101010101000010100001;
12'b100110100000: dataB <= 32'b00110001010111110100101011001000;
12'b100110100001: dataB <= 32'b00000111010011011000111001001001;
12'b100110100010: dataB <= 32'b00010011000111000101000110100011;
12'b100110100011: dataB <= 32'b00001011110000111101000010010111;
12'b100110100100: dataB <= 32'b01101100110010001011000111000111;
12'b100110100101: dataB <= 32'b00000110100001100000000111001100;
12'b100110100110: dataB <= 32'b01100101010011100100101111001101;
12'b100110100111: dataB <= 32'b00000000101100011111000000011010;
12'b100110101000: dataB <= 32'b00010100011110101011011010100111;
12'b100110101001: dataB <= 32'b00000111100011110100100011000111;
12'b100110101010: dataB <= 32'b01100100001101111001111000100001;
12'b100110101011: dataB <= 32'b00000110011000010010110101101000;
12'b100110101100: dataB <= 32'b11111001000101011100100010001000;
12'b100110101101: dataB <= 32'b00000011101010100011001010100011;
12'b100110101110: dataB <= 32'b00011010000101110111100000101011;
12'b100110101111: dataB <= 32'b00001001010111011111001010001010;
12'b100110110000: dataB <= 32'b11010000010111000101010110000111;
12'b100110110001: dataB <= 32'b00001010010001011010100010011100;
12'b100110110010: dataB <= 32'b10011011000100001011010010101100;
12'b100110110011: dataB <= 32'b00000011111100001101011010011111;
12'b100110110100: dataB <= 32'b01111100110110110010111001100101;
12'b100110110101: dataB <= 32'b00001000000001111101001011001010;
12'b100110110110: dataB <= 32'b01101100001110010010011110010000;
12'b100110110111: dataB <= 32'b00001000011100001100110010100010;
12'b100110111000: dataB <= 32'b01011011000100001100100010110100;
12'b100110111001: dataB <= 32'b00001011010111100111001010000101;
12'b100110111010: dataB <= 32'b10010001000100101100010111111100;
12'b100110111011: dataB <= 32'b00001110110000110100110000010010;
12'b100110111100: dataB <= 32'b00000000000001001001110110001010;
12'b100110111101: dataB <= 32'b00000000000000000000000000000000;
12'b100110111110: dataB <= 32'b10010000010100001011000001100111;
12'b100110111111: dataB <= 32'b00001000110101010110101010101111;
12'b100111000000: dataB <= 32'b00101110001101010111010100111000;
12'b100111000001: dataB <= 32'b00001110010111111011000010010001;
12'b100111000010: dataB <= 32'b10000011000111000100011011101011;
12'b100111000011: dataB <= 32'b00001100011100101011001100010101;
12'b100111000100: dataB <= 32'b10010100101100101100100101001111;
12'b100111000101: dataB <= 32'b00001010001011100110011010001111;
12'b100111000110: dataB <= 32'b10100010000110101101001010001111;
12'b100111000111: dataB <= 32'b00000011101100001010010111010101;
12'b100111001000: dataB <= 32'b01011011000010011111100111111000;
12'b100111001001: dataB <= 32'b00001010110101011000000101110101;
12'b100111001010: dataB <= 32'b01100010110010111011011101001000;
12'b100111001011: dataB <= 32'b00000111100110110011010110011100;
12'b100111001100: dataB <= 32'b11010101101011001010101100000100;
12'b100111001101: dataB <= 32'b00001101111001100110101000011101;
12'b100111001110: dataB <= 32'b10011101100001101110100111010100;
12'b100111001111: dataB <= 32'b00000100000011101001010100011011;
12'b100111010000: dataB <= 32'b01111000110011110101001100000011;
12'b100111010001: dataB <= 32'b00001011010100111001100011101100;
12'b100111010010: dataB <= 32'b00010000100011000100011111001101;
12'b100111010011: dataB <= 32'b00001010110010100100011000011010;
12'b100111010100: dataB <= 32'b00010100111101111011111001110100;
12'b100111010101: dataB <= 32'b00001101011010011010001001100101;
12'b100111010110: dataB <= 32'b01100000000101011111101000011110;
12'b100111010111: dataB <= 32'b00001010010010101111011010111100;
12'b100111011000: dataB <= 32'b00001100110001110010011010110100;
12'b100111011001: dataB <= 32'b00001001000001110000001100001100;
12'b100111011010: dataB <= 32'b10010101010010011110000101000100;
12'b100111011011: dataB <= 32'b00001010011110011100111100110011;
12'b100111011100: dataB <= 32'b00000011001001110111100110111001;
12'b100111011101: dataB <= 32'b00000111111101011001010101000111;
12'b100111011110: dataB <= 32'b11000110100000001011001000110110;
12'b100111011111: dataB <= 32'b00001101010100110000111101000101;
12'b100111100000: dataB <= 32'b01011001010101100011110111110011;
12'b100111100001: dataB <= 32'b00000010101100010110111000110101;
12'b100111100010: dataB <= 32'b11110110111111001110111000000110;
12'b100111100011: dataB <= 32'b00000000110001010001001010111010;
12'b100111100100: dataB <= 32'b11100000011011000111001000101111;
12'b100111100101: dataB <= 32'b00000111011110001100111010101011;
12'b100111100110: dataB <= 32'b10010110100110111010111001000010;
12'b100111100111: dataB <= 32'b00000100010101001110111101110011;
12'b100111101000: dataB <= 32'b11011011011010000111101000010111;
12'b100111101001: dataB <= 32'b00001001010111011100110001010110;
12'b100111101010: dataB <= 32'b11011111010100101010111000011100;
12'b100111101011: dataB <= 32'b00001101110100110010011000110010;
12'b100111101100: dataB <= 32'b11111100111111011110011100110001;
12'b100111101101: dataB <= 32'b00001001011010010100011110011010;
12'b100111101110: dataB <= 32'b10011001001001101010100101100011;
12'b100111101111: dataB <= 32'b00001000001010100000010001001101;
12'b100111110000: dataB <= 32'b01010101010010101001111111010001;
12'b100111110001: dataB <= 32'b00000110011000001100110001011110;
12'b100111110010: dataB <= 32'b01001001000010001110011000010100;
12'b100111110011: dataB <= 32'b00001100010011100100100000100110;
12'b100111110100: dataB <= 32'b10110010101010001001001010100001;
12'b100111110101: dataB <= 32'b00000101011100010100111110110001;
12'b100111110110: dataB <= 32'b11101101011011110101001011101001;
12'b100111110111: dataB <= 32'b00000111010011011000111001011000;
12'b100111111000: dataB <= 32'b00010011000010111101101000000011;
12'b100111111001: dataB <= 32'b00001011010010111101001101111111;
12'b100111111010: dataB <= 32'b11101100110110001011000111100111;
12'b100111111011: dataB <= 32'b00001000000001100110000111000100;
12'b100111111100: dataB <= 32'b10100011010011011101011111010000;
12'b100111111101: dataB <= 32'b00000001001001011111000000101001;
12'b100111111110: dataB <= 32'b01011000011010110011101011001001;
12'b100111111111: dataB <= 32'b00001001000011110110101010110111;
12'b101000000000: dataB <= 32'b01101010010010001001111010000010;
12'b101000000001: dataB <= 32'b00000101111000010010110010000000;
12'b101000000010: dataB <= 32'b00111001001101011100010011000110;
12'b101000000011: dataB <= 32'b00000100101001100011001010100100;
12'b101000000100: dataB <= 32'b00011110000101011111100001101000;
12'b101000000101: dataB <= 32'b00001000010111011111001010010010;
12'b101000000110: dataB <= 32'b11010100010010110101100111000110;
12'b101000000111: dataB <= 32'b00001010010010011110100010011100;
12'b101000001000: dataB <= 32'b10011001000000010010100011001010;
12'b101000001001: dataB <= 32'b00000010111010001011010010000111;
12'b101000001010: dataB <= 32'b11111101000010111011011010100101;
12'b101000001011: dataB <= 32'b00001001100001111101010111010010;
12'b101000001100: dataB <= 32'b10110000010010011010101101110010;
12'b101000001101: dataB <= 32'b00000110111100001110101010110010;
12'b101000001110: dataB <= 32'b01011011000100001100000010010010;
12'b101000001111: dataB <= 32'b00001010011000100101001101111101;
12'b101000010000: dataB <= 32'b11001110111100101011100110111011;
12'b101000010001: dataB <= 32'b00001110110011110100111000011001;
12'b101000010010: dataB <= 32'b00000000000001010001100111001010;
12'b101000010011: dataB <= 32'b00000000000000000000000000000000;
12'b101000010100: dataB <= 32'b10010100010000010010010010100100;
12'b101000010101: dataB <= 32'b00001000010110011010100110010111;
12'b101000010110: dataB <= 32'b01110010010001000110110011110110;
12'b101000010111: dataB <= 32'b00001101111010111001001110101001;
12'b101000011000: dataB <= 32'b11000010111011000100101100001101;
12'b101000011001: dataB <= 32'b00001011011101101001010000001100;
12'b101000011010: dataB <= 32'b10010110101000101100000101001110;
12'b101000011011: dataB <= 32'b00001010101100101010011001110111;
12'b101000011100: dataB <= 32'b00101000000110100101011010010000;
12'b101000011101: dataB <= 32'b00000100001011001110001111000110;
12'b101000011110: dataB <= 32'b00011010111110000111100111010111;
12'b101000011111: dataB <= 32'b00001001110110011110000101101101;
12'b101000100000: dataB <= 32'b10100100110111000011111101101010;
12'b101000100001: dataB <= 32'b00001000100110110001011010010100;
12'b101000100010: dataB <= 32'b01010001100111010011001101000110;
12'b101000100011: dataB <= 32'b00001100111011101000101100001101;
12'b101000100100: dataB <= 32'b00011011100001011110010111010011;
12'b101000100101: dataB <= 32'b00000101000001100101011000100011;
12'b101000100110: dataB <= 32'b00111010111111101101111101000101;
12'b101000100111: dataB <= 32'b00001010110101110101101111100101;
12'b101000101000: dataB <= 32'b10010100011111000100101111010000;
12'b101000101001: dataB <= 32'b00001010110011101000011100100001;
12'b101000101010: dataB <= 32'b11010100111001111011111001010101;
12'b101000101011: dataB <= 32'b00001011111100100000001001011100;
12'b101000101100: dataB <= 32'b11100100000101000111010110111110;
12'b101000101101: dataB <= 32'b00001010010010101101011110111100;
12'b101000101110: dataB <= 32'b01001100101010000010011010010101;
12'b101000101111: dataB <= 32'b00001010000001110100010100001011;
12'b101000110000: dataB <= 32'b00010011001010001110000110100011;
12'b101000110001: dataB <= 32'b00001000111110011100111100110011;
12'b101000110010: dataB <= 32'b11000010111101011111100101111000;
12'b101000110011: dataB <= 32'b00000110011100010111010000101110;
12'b101000110100: dataB <= 32'b01001000010100010010010111110110;
12'b101000110101: dataB <= 32'b00001100110110110001000100111101;
12'b101000110110: dataB <= 32'b11010111010001100011100111010011;
12'b101000110111: dataB <= 32'b00000011001010011000111000101100;
12'b101000111000: dataB <= 32'b01110111000110111111011001000110;
12'b101000111001: dataB <= 32'b00000000101110010001000111000011;
12'b101000111010: dataB <= 32'b00100100011010110111011000101111;
12'b101000111011: dataB <= 32'b00000101111110001110110010101100;
12'b101000111100: dataB <= 32'b10011000100011000011011010100010;
12'b101000111101: dataB <= 32'b00000011110011010000111001110011;
12'b101000111110: dataB <= 32'b10011001011001101111100111110111;
12'b101000111111: dataB <= 32'b00001000011000011100110001000110;
12'b101001000000: dataB <= 32'b10011101010100110010010111011011;
12'b101001000001: dataB <= 32'b00001101010110110110100000111010;
12'b101001000010: dataB <= 32'b00111101000111001110111100010011;
12'b101001000011: dataB <= 32'b00001000011010011000011010100011;
12'b101001000100: dataB <= 32'b01011001001001110010100111000010;
12'b101001000101: dataB <= 32'b00001000101010100100010001000101;
12'b101001000110: dataB <= 32'b00010011001010111010001111010100;
12'b101001000111: dataB <= 32'b00000101110111001100101001010110;
12'b101001001000: dataB <= 32'b11001000111001111110010111110100;
12'b101001001001: dataB <= 32'b00001011110100101000100100010101;
12'b101001001010: dataB <= 32'b00110100110010100001011011100011;
12'b101001001011: dataB <= 32'b00000011111010010100111011000010;
12'b101001001100: dataB <= 32'b10101011011111100101111100001011;
12'b101001001101: dataB <= 32'b00000110110010011010110101110000;
12'b101001001110: dataB <= 32'b00010010111010110101111001000011;
12'b101001001111: dataB <= 32'b00001011010011111011010101101111;
12'b101001010000: dataB <= 32'b00101100111010010011011000100111;
12'b101001010001: dataB <= 32'b00001001100001101100001010111101;
12'b101001010010: dataB <= 32'b01100001010111010101111111010010;
12'b101001010011: dataB <= 32'b00000001100111011111000000111001;
12'b101001010100: dataB <= 32'b10011100011010110100001011101010;
12'b101001010101: dataB <= 32'b00001010000100111000110110011111;
12'b101001010110: dataB <= 32'b01101110010110010001111011000011;
12'b101001010111: dataB <= 32'b00000100110111010100101110011000;
12'b101001011000: dataB <= 32'b01110111010101010100000100000100;
12'b101001011001: dataB <= 32'b00000101001000100001001010100100;
12'b101001011010: dataB <= 32'b01100100000101000111010010000110;
12'b101001011011: dataB <= 32'b00000111110111011101001010100010;
12'b101001011100: dataB <= 32'b00011010001110101101111000000110;
12'b101001011101: dataB <= 32'b00001010010010100000100010010101;
12'b101001011110: dataB <= 32'b10011000111100011001110011101001;
12'b101001011111: dataB <= 32'b00000001110111001011001001101111;
12'b101001100000: dataB <= 32'b01111101001010111011101011100111;
12'b101001100001: dataB <= 32'b00001010100010111001011111010011;
12'b101001100010: dataB <= 32'b11110100011010100010111101010101;
12'b101001100011: dataB <= 32'b00000101111011010000100010111010;
12'b101001100100: dataB <= 32'b01011011000000001011010010010000;
12'b101001100101: dataB <= 32'b00001001011001100101001101110101;
12'b101001100110: dataB <= 32'b01010000111000101011000101011010;
12'b101001100111: dataB <= 32'b00001110010101110101000000101001;
12'b101001101000: dataB <= 32'b00000000000001100001010111101001;
12'b101001101001: dataB <= 32'b00000000000000000000000000000000;
12'b101001101010: dataB <= 32'b10011000001100011001110100000011;
12'b101001101011: dataB <= 32'b00000111110110011100100101111111;
12'b101001101100: dataB <= 32'b10110110011000101110100011010100;
12'b101001101101: dataB <= 32'b00001100011100110111010110111001;
12'b101001101110: dataB <= 32'b00000010101110111101001100001111;
12'b101001101111: dataB <= 32'b00001001111110100111010100001100;
12'b101001110000: dataB <= 32'b10011000100100101011010101001101;
12'b101001110001: dataB <= 32'b00001010101101101110100001011111;
12'b101001110010: dataB <= 32'b10101110001010011101101010010001;
12'b101001110011: dataB <= 32'b00000100101001010010001010111110;
12'b101001110100: dataB <= 32'b00011010111101101111100110010111;
12'b101001110101: dataB <= 32'b00001001010110100100000101100101;
12'b101001110110: dataB <= 32'b10100100110111000100011110001100;
12'b101001110111: dataB <= 32'b00001001100110101101100010010100;
12'b101001111000: dataB <= 32'b10001101011111010011101110001000;
12'b101001111001: dataB <= 32'b00001011011101101010110000001100;
12'b101001111010: dataB <= 32'b10010111011101001110000110110011;
12'b101001111011: dataB <= 32'b00000110100001100011011000101010;
12'b101001111100: dataB <= 32'b10111011000111011110011110000111;
12'b101001111101: dataB <= 32'b00001010010110101111110011011101;
12'b101001111110: dataB <= 32'b00011000011010111101001111010011;
12'b101001111111: dataB <= 32'b00001010010100101100100000110001;
12'b101010000000: dataB <= 32'b10010100110101111011111000110101;
12'b101010000001: dataB <= 32'b00001010111110100100001001011100;
12'b101010000010: dataB <= 32'b00101010001000110110110101111110;
12'b101010000011: dataB <= 32'b00001001110011101001100010110101;
12'b101010000100: dataB <= 32'b11010000100010001010011001110110;
12'b101010000101: dataB <= 32'b00001011100011111000011100001010;
12'b101010000110: dataB <= 32'b10010011000101111110010111100010;
12'b101010000111: dataB <= 32'b00000111011110011100111100111010;
12'b101010001000: dataB <= 32'b00000010110001000111010100110111;
12'b101010001001: dataB <= 32'b00000101011011010101001100011110;
12'b101010001010: dataB <= 32'b11001110001100011001110111010110;
12'b101010001011: dataB <= 32'b00001011111000110001001100110100;
12'b101010001100: dataB <= 32'b01010101001101100011100111010011;
12'b101010001101: dataB <= 32'b00000011101000011000110100101100;
12'b101010001110: dataB <= 32'b11110101001110100111101010000111;
12'b101010001111: dataB <= 32'b00000000101011001110111111000011;
12'b101010010000: dataB <= 32'b01101000011110011111101000101111;
12'b101010010001: dataB <= 32'b00000100011101010000101010101100;
12'b101010010010: dataB <= 32'b10011100100011000011111011100100;
12'b101010010011: dataB <= 32'b00000011110001010000110001110011;
12'b101010010100: dataB <= 32'b00010111010101011111100110110111;
12'b101010010101: dataB <= 32'b00000111011000011110110000110110;
12'b101010010110: dataB <= 32'b00011011010101000001110110011011;
12'b101010010111: dataB <= 32'b00001100011000111000101001001010;
12'b101010011000: dataB <= 32'b01111011010010110111011011110101;
12'b101010011001: dataB <= 32'b00000110111010011100011010100011;
12'b101010011010: dataB <= 32'b11011001000101111010101000000010;
12'b101010011011: dataB <= 32'b00001001001010101000010100111100;
12'b101010011100: dataB <= 32'b10010011000111000010101110110111;
12'b101010011101: dataB <= 32'b00000100110110010000100001000101;
12'b101010011110: dataB <= 32'b00001010110001101110010111010100;
12'b101010011111: dataB <= 32'b00001011010110101010101000001101;
12'b101010100000: dataB <= 32'b10110100111010110001101101000101;
12'b101010100001: dataB <= 32'b00000010111001010100110111001010;
12'b101010100010: dataB <= 32'b10100111100011011110011100101101;
12'b101010100011: dataB <= 32'b00000110110010011010110110000000;
12'b101010100100: dataB <= 32'b11010010110110100110001010000100;
12'b101010100101: dataB <= 32'b00001010110100111001100001011110;
12'b101010100110: dataB <= 32'b10101111000010010011011001100111;
12'b101010100111: dataB <= 32'b00001011000010110000001110110101;
12'b101010101000: dataB <= 32'b11011111010111000110011110110101;
12'b101010101001: dataB <= 32'b00000010100101011111000001001000;
12'b101010101010: dataB <= 32'b10100000010110110100011100001100;
12'b101010101011: dataB <= 32'b00001011000101111010111110000111;
12'b101010101100: dataB <= 32'b10110010011110100010001100000101;
12'b101010101101: dataB <= 32'b00000100010101010110101010110000;
12'b101010101110: dataB <= 32'b10110011100001010011110101000011;
12'b101010101111: dataB <= 32'b00000110000111100001001010100100;
12'b101010110000: dataB <= 32'b10101010001000110110110011000100;
12'b101010110001: dataB <= 32'b00000110110111011101001010101010;
12'b101010110010: dataB <= 32'b00011110001010011110001001000110;
12'b101010110011: dataB <= 32'b00001001110011100100100010001101;
12'b101010110100: dataB <= 32'b10011000111100101001010100100111;
12'b101010110101: dataB <= 32'b00000000110101001001000001011111;
12'b101010110110: dataB <= 32'b11111011010111000100001100101001;
12'b101010110111: dataB <= 32'b00001100000011110101101011011011;
12'b101010111000: dataB <= 32'b01111000100010101011001100110111;
12'b101010111001: dataB <= 32'b00000100111010010100011110111011;
12'b101010111010: dataB <= 32'b01011011000000010010100010001110;
12'b101010111011: dataB <= 32'b00001000011001100011001101101101;
12'b101010111100: dataB <= 32'b11010000110000110010100100011001;
12'b101010111101: dataB <= 32'b00001101010111110101001100111000;
12'b101010111110: dataB <= 32'b00000000000001110001011000001001;
12'b101010111111: dataB <= 32'b00000000000000000000000000000000;
endcase
end
assign doA = dataA;
assign doB = dataB;
endmodule
