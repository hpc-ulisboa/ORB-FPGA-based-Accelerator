module rams_sp_rom1_4_sec (clk, enA, enB, addrA, addrB, doA, doB);
input clk;
input enA, enB;
input [10:0] addrA, addrB;
output [31:0] doA, doB;
(*rom_style = "block" *) reg [1375:0] dataA, dataB;
always @(posedge clk)
begin
if (enA)
case(addrA)
11'b00000000000: dataA <= 32'b11000111010001000111010001111000;
11'b00000000001: dataA <= 32'b00001011001111010011001011110011;
11'b00000000010: dataA <= 32'b01001010010111010110011010111001;
11'b00000000011: dataA <= 32'b00001101100101101000001100101010;
11'b00000000100: dataA <= 32'b10011011111010011010000111000111;
11'b00000000101: dataA <= 32'b00001111001011101010101110001111;
11'b00000000110: dataA <= 32'b10010011010001111110100111010101;
11'b00000000111: dataA <= 32'b00000110001010001110100111110100;
11'b00000001000: dataA <= 32'b11000100101010110010111000101011;
11'b00000001001: dataA <= 32'b00000101010111000101011111001001;
11'b00000001010: dataA <= 32'b11011111001011110100001011110010;
11'b00000001011: dataA <= 32'b00001011001100000010111110100100;
11'b00000001100: dataA <= 32'b01011010110110000001110101100011;
11'b00000001101: dataA <= 32'b00000011001101101110100010010011;
11'b00000001110: dataA <= 32'b10110001100001101001010011100100;
11'b00000001111: dataA <= 32'b00001110000111010110101010011111;
11'b00000010000: dataA <= 32'b11101111001111001101011001110010;
11'b00000010001: dataA <= 32'b00000000110011101100110101011110;
11'b00000010010: dataA <= 32'b11100000001011000000110011000100;
11'b00000010011: dataA <= 32'b00001011001010111000011110101000;
11'b00000010100: dataA <= 32'b10001101010010011010001000100001;
11'b00000010101: dataA <= 32'b00001010001011001110101000101110;
11'b00000010110: dataA <= 32'b00011101010101111100001010101101;
11'b00000010111: dataA <= 32'b00001110101001000100111010010101;
11'b00000011000: dataA <= 32'b01000010101111100110001111010011;
11'b00000011001: dataA <= 32'b00001001101100110000101010011010;
11'b00000011010: dataA <= 32'b10010011100001001011111011001011;
11'b00000011011: dataA <= 32'b00000001001001001100010001100111;
11'b00000011100: dataA <= 32'b01100101011011001011110001110001;
11'b00000011101: dataA <= 32'b00001111010000011111000101011110;
11'b00000011110: dataA <= 32'b11011101111011101101011100010101;
11'b00000011111: dataA <= 32'b00001110010100101001010111010110;
11'b00000100000: dataA <= 32'b01001001101001000111011011010000;
11'b00000100001: dataA <= 32'b00001011100111100100011110100110;
11'b00000100010: dataA <= 32'b10101001010101110100111001110001;
11'b00000100011: dataA <= 32'b00000100111001011011001110010110;
11'b00000100100: dataA <= 32'b11100100010111101010100011101100;
11'b00000100101: dataA <= 32'b00000110111110100001100001110001;
11'b00000100110: dataA <= 32'b10001110110011110010110111101110;
11'b00000100111: dataA <= 32'b00001110110101010111100010000010;
11'b00000101000: dataA <= 32'b01010001001001110001110001101001;
11'b00000101001: dataA <= 32'b00001001011000011011011101110100;
11'b00000101010: dataA <= 32'b00101011001111110100111011110001;
11'b00000101011: dataA <= 32'b00001100010000011001000011001110;
11'b00000101100: dataA <= 32'b11101011000101000110001101110010;
11'b00000101101: dataA <= 32'b00001011100110010010010001001101;
11'b00000101110: dataA <= 32'b11100110001011100001111010000111;
11'b00000101111: dataA <= 32'b00001101010000001101001001101010;
11'b00000110000: dataA <= 32'b00100011001101010100010001010000;
11'b00000110001: dataA <= 32'b00000101001110001010110010100110;
11'b00000110010: dataA <= 32'b10100101011001001010001010100010;
11'b00000110011: dataA <= 32'b00001011110101010011100010111101;
11'b00000110100: dataA <= 32'b01011011101011001100011010010001;
11'b00000110101: dataA <= 32'b00001010101000010010101110101111;
11'b00000110110: dataA <= 32'b11011010010100101010100010000110;
11'b00000110111: dataA <= 32'b00001100111001011101010101001001;
11'b00000111000: dataA <= 32'b00110000101111000001000110000110;
11'b00000111001: dataA <= 32'b00001001010010011011001000010100;
11'b00000111010: dataA <= 32'b11011101011011000010100010001100;
11'b00000111011: dataA <= 32'b00001001101010101110001011011100;
11'b00000111100: dataA <= 32'b00011110100001101011010011101101;
11'b00000111101: dataA <= 32'b00000000101010000100100010101010;
11'b00000111110: dataA <= 32'b11101011000011000001101010000001;
11'b00000111111: dataA <= 32'b00000011011011100001000000100101;
11'b00001000000: dataA <= 32'b10001011000010000010010101100111;
11'b00001000001: dataA <= 32'b00000010001010011100001111110011;
11'b00001000010: dataA <= 32'b10001100011101000011000010001000;
11'b00001000011: dataA <= 32'b00001011010110010101010100001010;
11'b00001000100: dataA <= 32'b11101110010101111101010010010110;
11'b00001000101: dataA <= 32'b00000011110100100100111110010010;
11'b00001000110: dataA <= 32'b11000010101111100110000010111010;
11'b00001000111: dataA <= 32'b00001011110001100101000101001010;
11'b00001001000: dataA <= 32'b10000111000111000010110011001110;
11'b00001001001: dataA <= 32'b00001001101100010000111010100011;
11'b00001001010: dataA <= 32'b11011111001100110110110100010111;
11'b00001001011: dataA <= 32'b00001011011101100011101011110100;
11'b00001001100: dataA <= 32'b01101000000101111001110100000111;
11'b00001001101: dataA <= 32'b00000001001000110010010001110001;
11'b00001001110: dataA <= 32'b00001110010001011010101011000101;
11'b00001001111: dataA <= 32'b00001101110101010001011001100010;
11'b00001010000: dataA <= 32'b01100001001001011111100111111011;
11'b00001010001: dataA <= 32'b00001100101110100110111010101100;
11'b00001010010: dataA <= 32'b01011011011101011110011101010110;
11'b00001010011: dataA <= 32'b00001011000100100010010100100110;
11'b00001010100: dataA <= 32'b00000000000000101100100100110000;
11'b00001010101: dataA <= 32'b00000000000000000000000000000000;
11'b00001010110: dataA <= 32'b01001101100001110111100100011100;
11'b00001010111: dataA <= 32'b00001010101101010101010011101010;
11'b00001011000: dataA <= 32'b10000100100111101101001100010110;
11'b00001011001: dataA <= 32'b00001011000010011110001000100011;
11'b00001011010: dataA <= 32'b00100111111010000001110101001000;
11'b00001011011: dataA <= 32'b00001101100110100110101010111111;
11'b00001011100: dataA <= 32'b00010111011010011110011000010101;
11'b00001011101: dataA <= 32'b00000101101100001010110111110011;
11'b00001011110: dataA <= 32'b00000011000010100010010111101011;
11'b00001011111: dataA <= 32'b00000110111000001101101110101001;
11'b00001100000: dataA <= 32'b01100001001011110010111100001111;
11'b00001100001: dataA <= 32'b00001010001010000011010010101100;
11'b00001100010: dataA <= 32'b00011000111001101010000011100110;
11'b00001100011: dataA <= 32'b00000011010001101000011010001011;
11'b00001100100: dataA <= 32'b11110111010001001001100001101000;
11'b00001100101: dataA <= 32'b00001100000011010100110011001110;
11'b00001100110: dataA <= 32'b00110001000011010100011010010000;
11'b00001100111: dataA <= 32'b00000010011001101010101101111111;
11'b00001101000: dataA <= 32'b10010110001110010000010001001001;
11'b00001101001: dataA <= 32'b00001001101000101110001110000000;
11'b00001101010: dataA <= 32'b01010011100010000001110110000001;
11'b00001101011: dataA <= 32'b00001000101001001100111001001111;
11'b00001101100: dataA <= 32'b11100001010101111100001010001011;
11'b00001101101: dataA <= 32'b00001100100100000101001110100100;
11'b00001101110: dataA <= 32'b00000011000111110100101111001101;
11'b00001101111: dataA <= 32'b00001000101011101010011110000010;
11'b00001110000: dataA <= 32'b10011011101001001100011010001001;
11'b00001110001: dataA <= 32'b00000000101111000100100110010111;
11'b00001110010: dataA <= 32'b01101001010111000010110010010110;
11'b00001110011: dataA <= 32'b00001110101010011111000101111110;
11'b00001110100: dataA <= 32'b10100111111011110011111100110001;
11'b00001110101: dataA <= 32'b00001110101111101011001111101101;
11'b00001110110: dataA <= 32'b10010011110101110111101011001110;
11'b00001110111: dataA <= 32'b00001001100101011100011111000101;
11'b00001111000: dataA <= 32'b01101011001110000100111001101111;
11'b00001111001: dataA <= 32'b00000110111011011111010010110110;
11'b00001111010: dataA <= 32'b00011100010011010001010011010000;
11'b00001111011: dataA <= 32'b00001001111110100111011101010010;
11'b00001111100: dataA <= 32'b10001101000011011001100111001110;
11'b00001111101: dataA <= 32'b00001111001111011101100101110010;
11'b00001111110: dataA <= 32'b01010011010101010010000000101110;
11'b00001111111: dataA <= 32'b00001010110110100001100001110100;
11'b00010000000: dataA <= 32'b11101101000111110011011011101110;
11'b00010000001: dataA <= 32'b00001011101101011001001011100100;
11'b00010000010: dataA <= 32'b01101010111101100110101101101110;
11'b00010000011: dataA <= 32'b00001001100100001010011101100110;
11'b00010000100: dataA <= 32'b00011010000111000000111000100110;
11'b00010000101: dataA <= 32'b00001100101100010001011001011011;
11'b00010000110: dataA <= 32'b01100111001001011100110010010101;
11'b00010000111: dataA <= 32'b00000101010000001001000010111101;
11'b00010001000: dataA <= 32'b11101001010100110010111000000001;
11'b00010001001: dataA <= 32'b00001100010010011011101011001100;
11'b00010001010: dataA <= 32'b10100011101111001011011010001111;
11'b00010001011: dataA <= 32'b00001001000111010000110111010110;
11'b00010001100: dataA <= 32'b10010010011000100011110000101100;
11'b00010001101: dataA <= 32'b00001110010100100001010100110010;
11'b00010001110: dataA <= 32'b01101010100010011000010100001000;
11'b00010001111: dataA <= 32'b00001001110001011101001100100101;
11'b00010010000: dataA <= 32'b10100001011010101001110001110001;
11'b00010010001: dataA <= 32'b00001000101001100010000111100011;
11'b00010010010: dataA <= 32'b11011000100101100011100011110001;
11'b00010010011: dataA <= 32'b00000000110000000010111010010001;
11'b00010010100: dataA <= 32'b11101000111010011000110111000001;
11'b00010010101: dataA <= 32'b00000101111110100001000000111110;
11'b00010010110: dataA <= 32'b00001111010001110010010100001010;
11'b00010010111: dataA <= 32'b00000001101110010010010011100010;
11'b00010011000: dataA <= 32'b00000110110000111011110001001101;
11'b00010011001: dataA <= 32'b00001100010011011011011000001100;
11'b00010011010: dataA <= 32'b11100100001110001101000011111010;
11'b00010011011: dataA <= 32'b00000101010111100100111010000010;
11'b00010011100: dataA <= 32'b01000011000111110100100100111101;
11'b00010011101: dataA <= 32'b00001011101110100101000001000011;
11'b00010011110: dataA <= 32'b00001001011010101010000011010010;
11'b00010011111: dataA <= 32'b00001000101011010001000110011011;
11'b00010100000: dataA <= 32'b01100001001101011111100101111001;
11'b00010100001: dataA <= 32'b00001101111001101011100111110011;
11'b00010100010: dataA <= 32'b10011100000101100010000010101011;
11'b00010100011: dataA <= 32'b00000000101110100110000101010001;
11'b00010100100: dataA <= 32'b10000110100001010011001000100100;
11'b00010100101: dataA <= 32'b00001110010001010111100101001010;
11'b00010100110: dataA <= 32'b11100011001010001111101001111010;
11'b00010100111: dataA <= 32'b00001100001010100100110010101011;
11'b00010101000: dataA <= 32'b01100001100010000110101101110001;
11'b00010101001: dataA <= 32'b00001000100010011010010101000111;
11'b00010101010: dataA <= 32'b00000000000000110101100101010010;
11'b00010101011: dataA <= 32'b00000000000000000000000000000000;
11'b00010101100: dataA <= 32'b00010101101110011111100110111110;
11'b00010101101: dataA <= 32'b00001010001011011001011011001001;
11'b00010101110: dataA <= 32'b11000010111111110011101101010010;
11'b00010101111: dataA <= 32'b00001000000001010100010000100100;
11'b00010110000: dataA <= 32'b01110001110001100001110100001010;
11'b00010110001: dataA <= 32'b00001011000010100000100111011110;
11'b00010110010: dataA <= 32'b11011101011110110110001001010101;
11'b00010110011: dataA <= 32'b00000100101110001011000111100001;
11'b00010110100: dataA <= 32'b11000101010110001010000110101100;
11'b00010110101: dataA <= 32'b00001000111001011001111010001000;
11'b00010110110: dataA <= 32'b10100011000111011001101011101100;
11'b00010110111: dataA <= 32'b00001001001001001001100110101011;
11'b00010111000: dataA <= 32'b00011000111101010010010010001010;
11'b00010111001: dataA <= 32'b00000011110101100000010110000011;
11'b00010111010: dataA <= 32'b11111000111100110010010000101101;
11'b00010111011: dataA <= 32'b00001001100001010010111111100101;
11'b00010111100: dataA <= 32'b11110000110011010011011010001111;
11'b00010111101: dataA <= 32'b00000100011100100110100110100110;
11'b00010111110: dataA <= 32'b11001100011001101000010000101110;
11'b00010111111: dataA <= 32'b00001000000111100100000101011000;
11'b00011000000: dataA <= 32'b10011001100101100001110011000100;
11'b00011000001: dataA <= 32'b00000111101001001101000101111111;
11'b00011000010: dataA <= 32'b01100101010101111100001001001010;
11'b00011000011: dataA <= 32'b00001010000001001011100010101100;
11'b00011000100: dataA <= 32'b00000101011011110011011110001000;
11'b00011000101: dataA <= 32'b00000111101011100010011001101010;
11'b00011000110: dataA <= 32'b00100011101001011100111000101000;
11'b00011000111: dataA <= 32'b00000000110101000010111010111111;
11'b00011001000: dataA <= 32'b01101101001110101010010011111010;
11'b00011001001: dataA <= 32'b00001101000101100001000110011110;
11'b00011001010: dataA <= 32'b00110011101111101010101100101110;
11'b00011001011: dataA <= 32'b00001101101010101101000011110100;
11'b00011001100: dataA <= 32'b11011111111010011111101010001100;
11'b00011001101: dataA <= 32'b00000111100100010110100011001100;
11'b00011001110: dataA <= 32'b10101101000010001100111001101110;
11'b00011001111: dataA <= 32'b00001001011011100001010011001101;
11'b00011010000: dataA <= 32'b10010100011010101000100011110011;
11'b00011010001: dataA <= 32'b00001100011100101101010101000010;
11'b00011010010: dataA <= 32'b11001111001110110000100111001110;
11'b00011010011: dataA <= 32'b00001110101010100101100001100010;
11'b00011010100: dataA <= 32'b10011001011101000010100001010100;
11'b00011010101: dataA <= 32'b00001100010100100111011101111100;
11'b00011010110: dataA <= 32'b10101100111011100010001011001011;
11'b00011010111: dataA <= 32'b00001011001010011011001111100011;
11'b00011011000: dataA <= 32'b01101010110110000110111101001001;
11'b00011011001: dataA <= 32'b00000111000100000100110010000110;
11'b00011011010: dataA <= 32'b10010000001110011000010110100111;
11'b00011011011: dataA <= 32'b00001100001001010111100001010011;
11'b00011011100: dataA <= 32'b10100111000101100101000011111001;
11'b00011011101: dataA <= 32'b00000101010010001011010011001100;
11'b00011011110: dataA <= 32'b11101101001100101011110101000010;
11'b00011011111: dataA <= 32'b00001100101110100011101011001011;
11'b00011100000: dataA <= 32'b01101011100110111010101001101101;
11'b00011100001: dataA <= 32'b00000111000110010001000011101101;
11'b00011100010: dataA <= 32'b10001100100100101100110000110001;
11'b00011100011: dataA <= 32'b00001110101111100101010100100011;
11'b00011100100: dataA <= 32'b01100100011001101000010011001100;
11'b00011100101: dataA <= 32'b00001001110000011111001100111110;
11'b00011100110: dataA <= 32'b10100111010110001001100010010101;
11'b00011100111: dataA <= 32'b00000111001001010110000111011010;
11'b00011101000: dataA <= 32'b10010100101101100011110100010100;
11'b00011101001: dataA <= 32'b00000001010110000011001101110001;
11'b00011101010: dataA <= 32'b01100110110001110000110100100010;
11'b00011101011: dataA <= 32'b00001000011110100001000001100111;
11'b00011101100: dataA <= 32'b00010011011101100010110011001101;
11'b00011101101: dataA <= 32'b00000001110011001010011111001001;
11'b00011101110: dataA <= 32'b10000111000100111100110001010010;
11'b00011101111: dataA <= 32'b00001100110000011111011100010101;
11'b00011110000: dataA <= 32'b11011010001110011100110110011101;
11'b00011110001: dataA <= 32'b00000110111001100010110101110010;
11'b00011110010: dataA <= 32'b00000101011111110011010111111110;
11'b00011110011: dataA <= 32'b00001011001011100100111101000100;
11'b00011110100: dataA <= 32'b11001111101010010001100100010101;
11'b00011110101: dataA <= 32'b00000111101011010011010010001010;
11'b00011110110: dataA <= 32'b00100011001010001111100111111010;
11'b00011110111: dataA <= 32'b00001111010100110001011011100010;
11'b00011111000: dataA <= 32'b01010010001001001010100010001111;
11'b00011111001: dataA <= 32'b00000000110100011100000100111010;
11'b00011111010: dataA <= 32'b01000010110101001011110110000100;
11'b00011111011: dataA <= 32'b00001110001100011111101001000011;
11'b00011111100: dataA <= 32'b01100101000110111111011011111000;
11'b00011111101: dataA <= 32'b00001010100111100010110010101011;
11'b00011111110: dataA <= 32'b10100111011110100110011101101100;
11'b00011111111: dataA <= 32'b00000110000010010010011101110111;
11'b00100000000: dataA <= 32'b00000000000001001110010101110100;
11'b00100000001: dataA <= 32'b00000000000000000000000000000000;
11'b00100000010: dataA <= 32'b01011111110111001110111001111110;
11'b00100000011: dataA <= 32'b00001001001010011111011110100000;
11'b00100000100: dataA <= 32'b11000011010111100010011101001110;
11'b00100000101: dataA <= 32'b00000101000001001100011000110101;
11'b00100000110: dataA <= 32'b11111001100001010010010011101110;
11'b00100000111: dataA <= 32'b00001000000001011100100111110100;
11'b00100001000: dataA <= 32'b11100011011111001101001010010011;
11'b00100001001: dataA <= 32'b00000100110000001101010111000000;
11'b00100001010: dataA <= 32'b00001011101001110010000110001101;
11'b00100001011: dataA <= 32'b00001010011000100011111001100001;
11'b00100001100: dataA <= 32'b00100011000110110000101010101001;
11'b00100001101: dataA <= 32'b00000111101000010011110110100011;
11'b00100001110: dataA <= 32'b00011001000101000011000001001111;
11'b00100001111: dataA <= 32'b00000101011000010110011001110011;
11'b00100010000: dataA <= 32'b01110110101100101011010001010011;
11'b00100010001: dataA <= 32'b00000110100001010011000111110100;
11'b00100010010: dataA <= 32'b00101100101011000010011001101101;
11'b00100010011: dataA <= 32'b00000111011110100000100011000110;
11'b00100010100: dataA <= 32'b10000110101000111000110000110100;
11'b00100010101: dataA <= 32'b00000110101000011000000100110001;
11'b00100010110: dataA <= 32'b10100001101001010010010001001000;
11'b00100010111: dataA <= 32'b00000110101010001111010110101111;
11'b00100011000: dataA <= 32'b11101001001101111100001000001001;
11'b00100011001: dataA <= 32'b00000111100001010011101110101011;
11'b00100011010: dataA <= 32'b01001101101111100001111100000011;
11'b00100011011: dataA <= 32'b00000110101011011010011001011010;
11'b00100011100: dataA <= 32'b00101011100101100101010111001000;
11'b00100011101: dataA <= 32'b00000010011010000011010011100110;
11'b00100011110: dataA <= 32'b11101111000010010001110110011100;
11'b00100011111: dataA <= 32'b00001010100010100001000110110101;
11'b00100100000: dataA <= 32'b10111011011111010001011100001010;
11'b00100100001: dataA <= 32'b00001100100110101100111011110010;
11'b00100100010: dataA <= 32'b11101011111011001110111001101010;
11'b00100100011: dataA <= 32'b00000101000101010000101011010011;
11'b00100100100: dataA <= 32'b10101100111010010100101001001101;
11'b00100100101: dataA <= 32'b00001011011001100101001111010100;
11'b00100100110: dataA <= 32'b10001110100101111000010100110110;
11'b00100100111: dataA <= 32'b00001110011000101111001000111011;
11'b00100101000: dataA <= 32'b01010011011010000000010111001111;
11'b00100101001: dataA <= 32'b00001101000101101011011101011011;
11'b00100101010: dataA <= 32'b10011111100000111011100010111001;
11'b00100101011: dataA <= 32'b00001100110000101101010110000100;
11'b00100101100: dataA <= 32'b10101010110011000000111010001001;
11'b00100101101: dataA <= 32'b00001001101000011111001111011010;
11'b00100101110: dataA <= 32'b01100110101110101110101011100110;
11'b00100101111: dataA <= 32'b00000100100101000101000110100110;
11'b00100110000: dataA <= 32'b00001000011101101000010101001000;
11'b00100110001: dataA <= 32'b00001010000110011111101001010100;
11'b00100110010: dataA <= 32'b10101000111101110101010101111100;
11'b00100110011: dataA <= 32'b00000110010100010001100011001011;
11'b00100110100: dataA <= 32'b11101111000000110100110010100101;
11'b00100110101: dataA <= 32'b00001100001011101011100111001010;
11'b00100110110: dataA <= 32'b11110001011010100001111001001100;
11'b00100110111: dataA <= 32'b00000101100111010011001111110011;
11'b00100111000: dataA <= 32'b10001010110100111101110001010111;
11'b00100111001: dataA <= 32'b00001110001010101001001100101100;
11'b00100111010: dataA <= 32'b00011100011001000000110010110000;
11'b00100111011: dataA <= 32'b00001001101110100011001101011111;
11'b00100111100: dataA <= 32'b10101011010001101001100011111001;
11'b00100111101: dataA <= 32'b00000110001010001100010011000001;
11'b00100111110: dataA <= 32'b11010010110101100100010101010111;
11'b00100111111: dataA <= 32'b00000010111010001001100101011001;
11'b00101000000: dataA <= 32'b01100010101101010001000010000110;
11'b00101000001: dataA <= 32'b00001011011101100001000010010111;
11'b00101000010: dataA <= 32'b01011011100101010011000011010001;
11'b00101000011: dataA <= 32'b00000011011000000110110010011000;
11'b00101000100: dataA <= 32'b10001001010101001101010010010111;
11'b00101000101: dataA <= 32'b00001100001100100101011000101110;
11'b00101000110: dataA <= 32'b00010000010110100100011000111101;
11'b00101000111: dataA <= 32'b00001000111001100000110101100011;
11'b00101001000: dataA <= 32'b11001101101111100001111010111110;
11'b00101001001: dataA <= 32'b00001010001001100100111001001100;
11'b00101001010: dataA <= 32'b10011001110001110001100101111000;
11'b00101001011: dataA <= 32'b00000110101011010111011001111010;
11'b00101001100: dataA <= 32'b11100101000110111111011010011001;
11'b00101001101: dataA <= 32'b00001111001111110101001111000000;
11'b00101001110: dataA <= 32'b00001000011001000011010010110011;
11'b00101001111: dataA <= 32'b00000010011001010000001000101011;
11'b00101010000: dataA <= 32'b00000101001101001100010100000110;
11'b00101010001: dataA <= 32'b00001100100111100111100100111100;
11'b00101010010: dataA <= 32'b11100101000011011110011101010101;
11'b00101010011: dataA <= 32'b00001000100110011110101110011010;
11'b00101010100: dataA <= 32'b10101101010110111101111100101000;
11'b00101010101: dataA <= 32'b00000011100101001100101010100111;
11'b00101010110: dataA <= 32'b00000000000001101110100110110101;
11'b00101010111: dataA <= 32'b00000000000000000000000000000000;
11'b00101011000: dataA <= 32'b11111011000011011001101111001100;
11'b00101011001: dataA <= 32'b00000101001101101111000000001010;
11'b00101011010: dataA <= 32'b01101011111001001000110111000101;
11'b00101011011: dataA <= 32'b00000000110101001101100110111110;
11'b00101011100: dataA <= 32'b01110000001101001101010111011000;
11'b00101011101: dataA <= 32'b00000000101111010011000110011000;
11'b00101011110: dataA <= 32'b11101110111010100001101001101011;
11'b00101011111: dataA <= 32'b00001000010110101011100100011001;
11'b00101100000: dataA <= 32'b11110101101001000100010110110011;
11'b00101100001: dataA <= 32'b00001100001011111100111000100100;
11'b00101100010: dataA <= 32'b11100010111000010010010100101010;
11'b00101100011: dataA <= 32'b00000100010000111011011001100010;
11'b00101100100: dataA <= 32'b01100011001101100101110111111101;
11'b00101100101: dataA <= 32'b00001100010101001101010001100100;
11'b00101100110: dataA <= 32'b01010110010001101110101001111101;
11'b00101100111: dataA <= 32'b00000000110010100011011010001000;
11'b00101101000: dataA <= 32'b11010100100101001001110110101100;
11'b00101101001: dataA <= 32'b00001111010001010000111111000001;
11'b00101101010: dataA <= 32'b01010101110000011110001010011110;
11'b00101101011: dataA <= 32'b00000100010010000011001100110110;
11'b00101101100: dataA <= 32'b10110100111101001101010100011101;
11'b00101101101: dataA <= 32'b00000101010010101011100011110010;
11'b00101101110: dataA <= 32'b10100110101110000100000100101111;
11'b00101101111: dataA <= 32'b00000000110000110111011001111010;
11'b00101110000: dataA <= 32'b00110111100100111000110001100111;
11'b00101110001: dataA <= 32'b00000101110010001101001001001101;
11'b00101110010: dataA <= 32'b11110010101010101100110100010001;
11'b00101110011: dataA <= 32'b00001101011011101001111011000000;
11'b00101110100: dataA <= 32'b01100000100000111011011110010011;
11'b00101110101: dataA <= 32'b00000001001010100010111110111010;
11'b00101110110: dataA <= 32'b01101110001000101001010101000111;
11'b00101110111: dataA <= 32'b00000011000110011100100101010000;
11'b00101111000: dataA <= 32'b01111100101011011001100101001100;
11'b00101111001: dataA <= 32'b00000010110101010101011101111001;
11'b00101111010: dataA <= 32'b01011100100110010011010110101101;
11'b00101111011: dataA <= 32'b00001100101001100110110110010001;
11'b00101111100: dataA <= 32'b00010011100000001100001011010110;
11'b00101111101: dataA <= 32'b00001100000011100100100001110110;
11'b00101111110: dataA <= 32'b00101101011000001011110111110001;
11'b00101111111: dataA <= 32'b00000010100101101110101001101101;
11'b00110000000: dataA <= 32'b11110001000001110110001100111010;
11'b00110000001: dataA <= 32'b00001000000110101010100110010011;
11'b00110000010: dataA <= 32'b00011000101000011001110100101011;
11'b00110000011: dataA <= 32'b00000100001100100111000001010001;
11'b00110000100: dataA <= 32'b11010110110011010010100011001000;
11'b00110000101: dataA <= 32'b00000010110110100011110111001010;
11'b00110000110: dataA <= 32'b01001111101100001100100100010101;
11'b00110000111: dataA <= 32'b00000011001011110101000010000101;
11'b00110001000: dataA <= 32'b10011110101110101100011110010100;
11'b00110001001: dataA <= 32'b00001010010011110001011101110001;
11'b00110001010: dataA <= 32'b10100000100010011110010010111010;
11'b00110001011: dataA <= 32'b00000101100111110010101001011001;
11'b00110001100: dataA <= 32'b01101100011100111010110110001101;
11'b00110001101: dataA <= 32'b00000011110100100111011001111000;
11'b00110001110: dataA <= 32'b10011011101010111110001011111101;
11'b00110001111: dataA <= 32'b00000101000011100110101110010110;
11'b00110010000: dataA <= 32'b00001101000100011101111000011010;
11'b00110010001: dataA <= 32'b00000111001100100110111011100101;
11'b00110010010: dataA <= 32'b11101000101000110100101100111000;
11'b00110010011: dataA <= 32'b00000101010011001001100100110001;
11'b00110010100: dataA <= 32'b00011011011010001100111011110101;
11'b00110010101: dataA <= 32'b00001101011010110011101100111101;
11'b00110010110: dataA <= 32'b01010110111000100101010011011011;
11'b00110010111: dataA <= 32'b00001110101001100000111111101011;
11'b00110011000: dataA <= 32'b00110011001001100101011000111001;
11'b00110011001: dataA <= 32'b00001100011001011001110000001011;
11'b00110011010: dataA <= 32'b10101011101110101101101011111011;
11'b00110011011: dataA <= 32'b00000110000111101100110111010110;
11'b00110011100: dataA <= 32'b11001011011110001010111110101110;
11'b00110011101: dataA <= 32'b00001100101110011010111101100100;
11'b00110011110: dataA <= 32'b10110111100100111000111111001010;
11'b00110011111: dataA <= 32'b00000100101011011100110110011101;
11'b00110100000: dataA <= 32'b00111001001100110100011100010100;
11'b00110100001: dataA <= 32'b00000101110010101101010001010100;
11'b00110100010: dataA <= 32'b11100010110111101010001100101011;
11'b00110100011: dataA <= 32'b00000111100001100110010100011001;
11'b00110100100: dataA <= 32'b10001101101101101101111001111010;
11'b00110100101: dataA <= 32'b00001100111011000101011101100110;
11'b00110100110: dataA <= 32'b00100111110110001101100011010111;
11'b00110100111: dataA <= 32'b00000011100110110010110010000110;
11'b00110101000: dataA <= 32'b00100000110111001001001010100101;
11'b00110101001: dataA <= 32'b00000011001110010111000001011011;
11'b00110101010: dataA <= 32'b11101010100110111010000100000110;
11'b00110101011: dataA <= 32'b00000010111000010101100111110010;
11'b00110101100: dataA <= 32'b00000000000011010100101010110010;
11'b00110101101: dataA <= 32'b00000000000000000000000000000000;
11'b00110101110: dataA <= 32'b10110111010111110011001111010010;
11'b00110101111: dataA <= 32'b00000101101011101101001100100001;
11'b00110110000: dataA <= 32'b11011111111001110000011001000101;
11'b00110110001: dataA <= 32'b00000000101111001001010110011110;
11'b00110110010: dataA <= 32'b00111000011100111100110101010111;
11'b00110110011: dataA <= 32'b00000001001001010010111111001001;
11'b00110110100: dataA <= 32'b11101111000111000010011010101101;
11'b00110110101: dataA <= 32'b00000111010110100011101000111000;
11'b00110110110: dataA <= 32'b10101011110101000011100110010010;
11'b00110110111: dataA <= 32'b00001100101110111101001100011011;
11'b00110111000: dataA <= 32'b10100010111000110001000110001000;
11'b00110111001: dataA <= 32'b00000100101101110011101101110010;
11'b00110111010: dataA <= 32'b11011111001101001101010101011011;
11'b00110111011: dataA <= 32'b00001010111000001010111101100011;
11'b00110111100: dataA <= 32'b11011110001101001110010110111110;
11'b00110111101: dataA <= 32'b00000000101100011111011010111000;
11'b00110111110: dataA <= 32'b11011000011101101001010111101011;
11'b00110111111: dataA <= 32'b00001110010111010010110011011010;
11'b00111000000: dataA <= 32'b00001101100100001100100111011110;
11'b00111000001: dataA <= 32'b00000011101111000010110100011101;
11'b00111000010: dataA <= 32'b00110011001100111100110010011001;
11'b00111000011: dataA <= 32'b00000100110000100011100111110100;
11'b00111000100: dataA <= 32'b10101010110110000100000101001101;
11'b00111000101: dataA <= 32'b00000000101011110001101010001010;
11'b00111000110: dataA <= 32'b10101101110101101000010100000011;
11'b00111000111: dataA <= 32'b00000101110000001100111001000100;
11'b00111001000: dataA <= 32'b00110100111010011101000100001110;
11'b00111001001: dataA <= 32'b00001010111110011101111011100010;
11'b00111001010: dataA <= 32'b00100110100101001010101101011000;
11'b00111001011: dataA <= 32'b00000010100101100010111111001011;
11'b00111001100: dataA <= 32'b01110110011001010000100111000110;
11'b00111001101: dataA <= 32'b00000101000100100000100110000000;
11'b00111001110: dataA <= 32'b10111101000011110011000110001011;
11'b00111001111: dataA <= 32'b00000010010000010001010010011001;
11'b00111010000: dataA <= 32'b10100000100110011011100111001100;
11'b00111010001: dataA <= 32'b00001101101101101000111110110001;
11'b00111010010: dataA <= 32'b11001101010100010010101001111000;
11'b00111010011: dataA <= 32'b00001110000111101010100101010101;
11'b00111010100: dataA <= 32'b11100111100000010010010111010001;
11'b00111010101: dataA <= 32'b00000101000010110000110101011100;
11'b00111010110: dataA <= 32'b00101111001101010101111010011101;
11'b00111010111: dataA <= 32'b00001010000111101110110010010100;
11'b00111011000: dataA <= 32'b11011100100101000000110101101001;
11'b00111011001: dataA <= 32'b00000101001001100111001001110000;
11'b00111011010: dataA <= 32'b11011010101011011011110100100101;
11'b00111011011: dataA <= 32'b00000010010001011001110111001011;
11'b00111011100: dataA <= 32'b01000111011100001011000011110010;
11'b00111011101: dataA <= 32'b00000100100111110001010001110101;
11'b00111011110: dataA <= 32'b10100010110010100100111100111000;
11'b00111011111: dataA <= 32'b00001001010101101001101010010001;
11'b00111100000: dataA <= 32'b10100110100101111110100001010101;
11'b00111100001: dataA <= 32'b00000111000110110100111001111001;
11'b00111100010: dataA <= 32'b10110010101001010010000110101100;
11'b00111100011: dataA <= 32'b00000011010001100001011110101000;
11'b00111100100: dataA <= 32'b11010011100110011110101000111110;
11'b00111100101: dataA <= 32'b00000111100010101010110101110110;
11'b00111100110: dataA <= 32'b00001100110100001100100110011001;
11'b00111100111: dataA <= 32'b00001000001100100111000011001110;
11'b00111101000: dataA <= 32'b00101010110000110011101010111011;
11'b00111101001: dataA <= 32'b00000100110001000011010001010001;
11'b00111101010: dataA <= 32'b01010111010101111100111010010111;
11'b00111101011: dataA <= 32'b00001011011101100111111000110100;
11'b00111101100: dataA <= 32'b11011000110000011100010001010110;
11'b00111101101: dataA <= 32'b00001111001111100000111111101100;
11'b00111101110: dataA <= 32'b10101111011001011100110110111001;
11'b00111101111: dataA <= 32'b00001001111100001111101000100001;
11'b00111110000: dataA <= 32'b01100011110010011110001001011101;
11'b00111110001: dataA <= 32'b00001000000110101111000010110111;
11'b00111110010: dataA <= 32'b01000111001010011011001110110011;
11'b00111110011: dataA <= 32'b00001100110010011010111001011100;
11'b00111110100: dataA <= 32'b11101111110101101000011111010000;
11'b00111110101: dataA <= 32'b00000101101001011110110110000101;
11'b00111110110: dataA <= 32'b10110101100000110011011010110111;
11'b00111110111: dataA <= 32'b00000101110000101001011001011011;
11'b00111111000: dataA <= 32'b11100100111011110011101101010000;
11'b00111111001: dataA <= 32'b00001010000001101100011101000000;
11'b00111111010: dataA <= 32'b00000101011001010101100111111011;
11'b00111111011: dataA <= 32'b00001010011110000011000101001110;
11'b00111111100: dataA <= 32'b11011011111001111101100010010011;
11'b00111111101: dataA <= 32'b00000110000011110101000001101101;
11'b00111111110: dataA <= 32'b10100010110111101010001100001000;
11'b00111111111: dataA <= 32'b00000011101010011000111001101010;
11'b01000000000: dataA <= 32'b01101110110011001010110110000100;
11'b01000000001: dataA <= 32'b00000001010011001111011011110100;
11'b01000000010: dataA <= 32'b00000000000011001101101010010100;
11'b01000000011: dataA <= 32'b00000000000000000000000000000000;
11'b01000000100: dataA <= 32'b10110001100111110100011110010111;
11'b01000000101: dataA <= 32'b00000110101010101001010101001000;
11'b01000000110: dataA <= 32'b11010011110110100000101011000111;
11'b01000000111: dataA <= 32'b00000001001001000101000001110110;
11'b01000001000: dataA <= 32'b00111100110000111011110100010101;
11'b01000001001: dataA <= 32'b00000011000100010100110011100010;
11'b01000001010: dataA <= 32'b01101101010011001011001010101111;
11'b01000001011: dataA <= 32'b00000110010100011011101001100000;
11'b01000001100: dataA <= 32'b10100001111001001010110101110000;
11'b01000001101: dataA <= 32'b00001100010010110111100100100010;
11'b01000001110: dataA <= 32'b10100100111101011000010111100111;
11'b01000001111: dataA <= 32'b00000101001011101001111010001010;
11'b01000010000: dataA <= 32'b10011101001101000100100011011000;
11'b01000010001: dataA <= 32'b00001000111001001100101101100011;
11'b01000010010: dataA <= 32'b10101000010000110101100100011100;
11'b01000010011: dataA <= 32'b00000001100111011001010111011001;
11'b01000010100: dataA <= 32'b00100000011110001001011000001011;
11'b01000010101: dataA <= 32'b00001100111011010110101011100100;
11'b01000010110: dataA <= 32'b11000111010000001011010100111101;
11'b01000010111: dataA <= 32'b00000100001100000110100000010011;
11'b01000011000: dataA <= 32'b10110001011000111011110000110011;
11'b01000011001: dataA <= 32'b00000100101110011101100111101101;
11'b01000011010: dataA <= 32'b11101010111110000100000101101011;
11'b01000011011: dataA <= 32'b00000010000110100111110110011010;
11'b01000011100: dataA <= 32'b11100011111010010000010110100001;
11'b01000011101: dataA <= 32'b00000101101110001110101001000011;
11'b01000011110: dataA <= 32'b01110101001010001101100100101011;
11'b01000011111: dataA <= 32'b00000111111110010011110111110011;
11'b01000100000: dataA <= 32'b00101010101101011001111011011011;
11'b01000100001: dataA <= 32'b00000101000010100011000011001100;
11'b01000100010: dataA <= 32'b10111100110001111000011000100110;
11'b01000100011: dataA <= 32'b00000111100010100110101010110000;
11'b01000100100: dataA <= 32'b11111011011011110100010111001001;
11'b01000100101: dataA <= 32'b00000010101100001111000110110001;
11'b01000100110: dataA <= 32'b01100110101010011011110111101100;
11'b01000100111: dataA <= 32'b00001101110010101001000011001010;
11'b01000101000: dataA <= 32'b01001001000100101001011000011001;
11'b01000101001: dataA <= 32'b00001111001100101110110001000101;
11'b01000101010: dataA <= 32'b01100001100100110001000111010001;
11'b01000101011: dataA <= 32'b00000111100001110011000101010100;
11'b01000101100: dataA <= 32'b01101011011001000101010111011110;
11'b01000101101: dataA <= 32'b00001011001010110000111110001100;
11'b01000101110: dataA <= 32'b11100010100101101000010111001000;
11'b01000101111: dataA <= 32'b00000110101000100101001110011000;
11'b01000110000: dataA <= 32'b11011110101011010100110111000100;
11'b01000110001: dataA <= 32'b00000010001100001111101011001100;
11'b01000110010: dataA <= 32'b00000011001000011001110011001110;
11'b01000110011: dataA <= 32'b00000110000110101101011101100101;
11'b01000110100: dataA <= 32'b00100100110010011101001010111011;
11'b01000110101: dataA <= 32'b00001000010101100001101110101010;
11'b01000110110: dataA <= 32'b10101010101101011110010000101111;
11'b01000110111: dataA <= 32'b00001001000111110101001010011001;
11'b01000111000: dataA <= 32'b01110110111001101001100111101011;
11'b01000111001: dataA <= 32'b00000011101101011011011111010001;
11'b01000111010: dataA <= 32'b01001101011001111110110110011110;
11'b01000111011: dataA <= 32'b00001010000011101010111101010110;
11'b01000111100: dataA <= 32'b11010000101000001011000100010111;
11'b01000111101: dataA <= 32'b00001000101100100111000110101110;
11'b01000111110: dataA <= 32'b11101100111100111010101000111100;
11'b01000111111: dataA <= 32'b00000100101110000010111001110000;
11'b01001000000: dataA <= 32'b01010011001101110100111000111000;
11'b01001000001: dataA <= 32'b00001000011110011101111000111011;
11'b01001000010: dataA <= 32'b00011100101100011011000000110001;
11'b01001000011: dataA <= 32'b00001111010100100000111111011110;
11'b01001000100: dataA <= 32'b11101001100001001100010101010111;
11'b01001000101: dataA <= 32'b00000111011100001001011001000000;
11'b01001000110: dataA <= 32'b10011001110001111110000110111101;
11'b01001000111: dataA <= 32'b00001001100111101101001010000111;
11'b01001001000: dataA <= 32'b11000110110110100011101101011000;
11'b01001001001: dataA <= 32'b00001011110101011100110101011011;
11'b01001001010: dataA <= 32'b11100011111010010000011110110110;
11'b01001001011: dataA <= 32'b00000111001000100000110101101101;
11'b01001001100: dataA <= 32'b00101101101101000010101001011001;
11'b01001001101: dataA <= 32'b00000101101110100011011101100011;
11'b01001001110: dataA <= 32'b01100110111111110101001100110100;
11'b01001001111: dataA <= 32'b00001100100100110010101001101000;
11'b01001010000: dataA <= 32'b01000011000101000100110101111010;
11'b01001010001: dataA <= 32'b00000111011110000010110000110101;
11'b01001010010: dataA <= 32'b10010001110001100101010010001110;
11'b01001010011: dataA <= 32'b00001000100011110011010001010101;
11'b01001010100: dataA <= 32'b10100100111011110011101101001100;
11'b01001010101: dataA <= 32'b00000101000111011000110101111010;
11'b01001010110: dataA <= 32'b11110000111111010011111000100100;
11'b01001010111: dataA <= 32'b00000001001110001011001011101101;
11'b01001011000: dataA <= 32'b00000000000010110110011001010101;
11'b01001011001: dataA <= 32'b00000000000000000000000000000000;
11'b01001011010: dataA <= 32'b01101001110011101101111100011100;
11'b01001011011: dataA <= 32'b00000111101001100101011001111000;
11'b01001011100: dataA <= 32'b10001011101011001001011100101010;
11'b01001011101: dataA <= 32'b00000010100100000110101101001110;
11'b01001011110: dataA <= 32'b10111101001001000011000011110001;
11'b01001011111: dataA <= 32'b00000101100001010110101011110011;
11'b01001100000: dataA <= 32'b01101001011011010100001010110001;
11'b01001100001: dataA <= 32'b00000101010011010011100010010000;
11'b01001100010: dataA <= 32'b10010101110101011010010101101110;
11'b01001100011: dataA <= 32'b00001011110101101111110100111001;
11'b01001100100: dataA <= 32'b11100101000010000000011001001000;
11'b01001100101: dataA <= 32'b00000110001001011111111010011010;
11'b01001100110: dataA <= 32'b01011011001000111011110001110100;
11'b01001100111: dataA <= 32'b00000110111001010000100001101011;
11'b01001101000: dataA <= 32'b00110000011100101100100010011000;
11'b01001101001: dataA <= 32'b00000011100011010101010011110011;
11'b01001101010: dataA <= 32'b00100110100010101001101001001100;
11'b01001101011: dataA <= 32'b00001001111110011010100111011101;
11'b01001101100: dataA <= 32'b10000100111100011001110010011001;
11'b01001101101: dataA <= 32'b00000101001001001110001100011010;
11'b01001101110: dataA <= 32'b10101001100101000011000000101110;
11'b01001101111: dataA <= 32'b00000101101011010101100011010110;
11'b01001110000: dataA <= 32'b01101011000110000100000110101010;
11'b01001110001: dataA <= 32'b00000100100010011101110110100011;
11'b01001110010: dataA <= 32'b00010111111011000000111001100001;
11'b01001110011: dataA <= 32'b00000110001100010100011101001011;
11'b01001110100: dataA <= 32'b11110001011001111101100101101001;
11'b01001110101: dataA <= 32'b00000100111101001001100111110100;
11'b01001110110: dataA <= 32'b00101100110101111001101000111100;
11'b01001110111: dataA <= 32'b00001000000001100011000011001101;
11'b01001111000: dataA <= 32'b01111101000110101000101010100111;
11'b01001111001: dataA <= 32'b00001010000011101010101111011001;
11'b01001111010: dataA <= 32'b11110101101111101101111000001001;
11'b01001111011: dataA <= 32'b00000011101000001110110111001010;
11'b01001111100: dataA <= 32'b01101010101110011100011000101100;
11'b01001111101: dataA <= 32'b00001100110110100111001011010011;
11'b01001111110: dataA <= 32'b01001010110101010000100110011000;
11'b01001111111: dataA <= 32'b00001111010010110000111100111100;
11'b01010000000: dataA <= 32'b11011001100001011000010111010000;
11'b01010000001: dataA <= 32'b00001010100010110001010001010011;
11'b01010000010: dataA <= 32'b01100101011100111100010100111100;
11'b01010000011: dataA <= 32'b00001100001101101111001010001100;
11'b01010000100: dataA <= 32'b10100110101010011000011000101000;
11'b01010000101: dataA <= 32'b00001000000111100001001111000001;
11'b01010000110: dataA <= 32'b10100010101011000101111001000100;
11'b01010000111: dataA <= 32'b00000011001000001001011010111101;
11'b01010001000: dataA <= 32'b10000100110000111000110011101011;
11'b01010001001: dataA <= 32'b00001000000101100101100101011100;
11'b01010001010: dataA <= 32'b11100110111010001101011000011101;
11'b01010001011: dataA <= 32'b00000111010101011001101011000010;
11'b01010001100: dataA <= 32'b00101100110101000101100001001010;
11'b01010001101: dataA <= 32'b00001010101000110001011010110010;
11'b01010001110: dataA <= 32'b10110101001010001001101000101011;
11'b01010001111: dataA <= 32'b00000100001010010111011011101010;
11'b01010010000: dataA <= 32'b10001011001001010110100011011011;
11'b01010010001: dataA <= 32'b00001100100110101011000100111101;
11'b01010010010: dataA <= 32'b01010110011100100001110011010011;
11'b01010010011: dataA <= 32'b00001001001101100101001010000111;
11'b01010010100: dataA <= 32'b00101101000101010001110110011011;
11'b01010010101: dataA <= 32'b00000101001100000100100010011001;
11'b01010010110: dataA <= 32'b10010001000001101100100110111000;
11'b01010010111: dataA <= 32'b00000101011110010001110101000010;
11'b01010011000: dataA <= 32'b11100000101000110001110000101011;
11'b01010011001: dataA <= 32'b00001101111001100000111110111110;
11'b01010011010: dataA <= 32'b01100001101001001011110011110100;
11'b01010011011: dataA <= 32'b00000101011011000111000101110000;
11'b01010011100: dataA <= 32'b10001111100101100101110100011011;
11'b01010011101: dataA <= 32'b00001011001001101011010101010111;
11'b01010011110: dataA <= 32'b01001010100010101100001011011011;
11'b01010011111: dataA <= 32'b00001010011000011110110101011011;
11'b01010100000: dataA <= 32'b10010111111011000000111101011010;
11'b01010100001: dataA <= 32'b00001000101000100010110101011101;
11'b01010100010: dataA <= 32'b11100011110001011001110111011001;
11'b01010100011: dataA <= 32'b00000110001100011101011101110010;
11'b01010100100: dataA <= 32'b01100111000011011110011011110111;
11'b01010100101: dataA <= 32'b00001110101001110100111010011000;
11'b01010100110: dataA <= 32'b01000010101100111100000011110111;
11'b01010100111: dataA <= 32'b00000100011101001000011000101100;
11'b01010101000: dataA <= 32'b11001001100001010101000010101001;
11'b01010101001: dataA <= 32'b00001010100100101101011101000100;
11'b01010101010: dataA <= 32'b10100100111111110101001101110000;
11'b01010101011: dataA <= 32'b00000111000110011100110010001010;
11'b01010101100: dataA <= 32'b11101111001011001101001011000101;
11'b01010101101: dataA <= 32'b00000010001001001010111011001110;
11'b01010101110: dataA <= 32'b00000000000010010110101000010110;
11'b01010101111: dataA <= 32'b00000000000000000000000000000000;
11'b01010110000: dataA <= 32'b00111000101110111000101110000111;
11'b01010110001: dataA <= 32'b00000100110000101100110100001100;
11'b01010110010: dataA <= 32'b10110101101000101001100101000110;
11'b01010110011: dataA <= 32'b00000010011010010111110011010101;
11'b01010110100: dataA <= 32'b01100100000101100101111000111000;
11'b01010110101: dataA <= 32'b00000000110100010101010001110000;
11'b01010110110: dataA <= 32'b01101100101110000001011000101010;
11'b01010110111: dataA <= 32'b00001001110101110001011000001011;
11'b01010111000: dataA <= 32'b00111011010101001101000111010100;
11'b01010111001: dataA <= 32'b00001010101000111010100000110110;
11'b01010111010: dataA <= 32'b00100000110100001011110100001101;
11'b01010111011: dataA <= 32'b00000100110011111101000001011011;
11'b01010111100: dataA <= 32'b10100101001001111110001010011100;
11'b01010111101: dataA <= 32'b00001100110010010001011101101100;
11'b01010111110: dataA <= 32'b01001110011110010110101100011011;
11'b01010111111: dataA <= 32'b00000001111000101001010101100000;
11'b01011000000: dataA <= 32'b00010000110000110010100110001101;
11'b01011000001: dataA <= 32'b00001111001100010011001010100001;
11'b01011000010: dataA <= 32'b00011111110100111111001100111011;
11'b01011000011: dataA <= 32'b00000100110101000111100001010111;
11'b01011000100: dataA <= 32'b01110010101101100101110111011110;
11'b01011000101: dataA <= 32'b00000101110100110001010111010001;
11'b01011000110: dataA <= 32'b11100010101010000011110101010010;
11'b01011000111: dataA <= 32'b00000001010110111011000101101010;
11'b01011001000: dataA <= 32'b10111101010000011001110000101100;
11'b01011001001: dataA <= 32'b00000110010011001111010101100101;
11'b01011001010: dataA <= 32'b01101100011110110100000100110100;
11'b01011001011: dataA <= 32'b00001110110110110011101110011000;
11'b01011001100: dataA <= 32'b10011010100100110100001110001110;
11'b01011001101: dataA <= 32'b00000000101111100000111010100001;
11'b01011001110: dataA <= 32'b00100010000100010010100011101010;
11'b01011001111: dataA <= 32'b00000001101011010110101000101001;
11'b01011010000: dataA <= 32'b10110110010110111000100100101111;
11'b01011010001: dataA <= 32'b00000100011000011011100001011001;
11'b01011010010: dataA <= 32'b01010110101010001011000110001110;
11'b01011010011: dataA <= 32'b00001011000110100100110001101001;
11'b01011010100: dataA <= 32'b00011011101000010101011100010011;
11'b01011010101: dataA <= 32'b00001001000001011110011110001110;
11'b01011010110: dataA <= 32'b01110001001100001101001000010001;
11'b01011010111: dataA <= 32'b00000001001010101000011101111101;
11'b01011011000: dataA <= 32'b10101110110110001110001110010110;
11'b01011011001: dataA <= 32'b00000110100111100100100010001011;
11'b01011011010: dataA <= 32'b11010100110000001011000100001110;
11'b01011011011: dataA <= 32'b00000011101111100110111100110001;
11'b01011011100: dataA <= 32'b00010100111010111001110010001101;
11'b01011011101: dataA <= 32'b00000100011001101101101110110010;
11'b01011011110: dataA <= 32'b00011001110100011110000101111000;
11'b01011011111: dataA <= 32'b00000010101111110010110110010101;
11'b01011100000: dataA <= 32'b11011100110010101011101110101111;
11'b01011100001: dataA <= 32'b00001010110001110101001101011001;
11'b01011100010: dataA <= 32'b01011010100110110101110101011101;
11'b01011100011: dataA <= 32'b00000100001010101100011101000010;
11'b01011100100: dataA <= 32'b10100100010100110011100101101110;
11'b01011100101: dataA <= 32'b00000101010111101101010001010000;
11'b01011100110: dataA <= 32'b00100101101011010101011101111001;
11'b01011100111: dataA <= 32'b00000011000110100010101010110110;
11'b01011101000: dataA <= 32'b11001111010000111110111001111001;
11'b01011101001: dataA <= 32'b00000110101101100100110111101011;
11'b01011101010: dataA <= 32'b00100010100100111101011101110011;
11'b01011101011: dataA <= 32'b00000110010101010001110100100011;
11'b01011101100: dataA <= 32'b11100001011110010100101100010010;
11'b01011101101: dataA <= 32'b00001111010101111011011101010101;
11'b01011101110: dataA <= 32'b00010100111100111110010101111110;
11'b01011101111: dataA <= 32'b00001100100100011110111111011010;
11'b01011110000: dataA <= 32'b01110100111101111101101010011000;
11'b01011110001: dataA <= 32'b00001101110101100011110000001100;
11'b01011110010: dataA <= 32'b01110011100010111100111101110111;
11'b01011110011: dataA <= 32'b00000100101001101010101011110101;
11'b01011110100: dataA <= 32'b00010001101010000010101101101001;
11'b01011110101: dataA <= 32'b00001100001011011011000001101101;
11'b01011110110: dataA <= 32'b00111101010000011001111101000101;
11'b01011110111: dataA <= 32'b00000100001110011010111010110101;
11'b01011111000: dataA <= 32'b01111000111000111101001100110001;
11'b01011111001: dataA <= 32'b00000110010011101111000101011100;
11'b01011111010: dataA <= 32'b00100000110011001001001011101000;
11'b01011111011: dataA <= 32'b00000100100010011100010100001011;
11'b01011111100: dataA <= 32'b10010111111010000110001011111000;
11'b01011111101: dataA <= 32'b00001110110111001101101110001110;
11'b01011111110: dataA <= 32'b11110001101110100101010100111010;
11'b01011111111: dataA <= 32'b00000010001010101110100110011101;
11'b01100000000: dataA <= 32'b10011110110110100000011000000100;
11'b01100000001: dataA <= 32'b00000011010001011001000101010011;
11'b01100000010: dataA <= 32'b10100100100010100001100010101001;
11'b01100000011: dataA <= 32'b00000100111011011101101011011001;
11'b01100000100: dataA <= 32'b00000000000011010011011011001111;
11'b01100000101: dataA <= 32'b00000000000000000000000000000000;
11'b01100000110: dataA <= 32'b10110010011110001000011011100011;
11'b01100000111: dataA <= 32'b00000101010010101010101100010101;
11'b01100001000: dataA <= 32'b01111011011000010010110011101001;
11'b01100001001: dataA <= 32'b00000100111101100001110111011100;
11'b01100001010: dataA <= 32'b11011000000101111110001010110111;
11'b01100001011: dataA <= 32'b00000010011001011001010101000000;
11'b01100001100: dataA <= 32'b11101000100101100001100111101010;
11'b01100001101: dataA <= 32'b00001010010011110101001000001100;
11'b01100001110: dataA <= 32'b11111100111101011101101000010100;
11'b01100001111: dataA <= 32'b00001001000111110010010001010110;
11'b01100010000: dataA <= 32'b10011110110100001101000011110000;
11'b01100010001: dataA <= 32'b00000101110101111100101101010011;
11'b01100010010: dataA <= 32'b11100111000110010101111100011001;
11'b01100010011: dataA <= 32'b00001100101110010111100101110100;
11'b01100010100: dataA <= 32'b00001000101110110110011110010111;
11'b01100010101: dataA <= 32'b00000011111100101011001100110001;
11'b01100010110: dataA <= 32'b11001110111100101011100101101111;
11'b01100010111: dataA <= 32'b00001101100110010101010010000000;
11'b01100011000: dataA <= 32'b01101001110001101111101110110110;
11'b01100011001: dataA <= 32'b00000110010111010001110001111111;
11'b01100011010: dataA <= 32'b10101100011101111110001001111110;
11'b01100011011: dataA <= 32'b00000111010110110011000110110000;
11'b01100011100: dataA <= 32'b00011110101010000011110101110100;
11'b01100011101: dataA <= 32'b00000011011011111010110001011011;
11'b01100011110: dataA <= 32'b11111100111000001011010000110010;
11'b01100011111: dataA <= 32'b00000111010100010101100001111101;
11'b01100100000: dataA <= 32'b01100100010110110011100101110110;
11'b01100100001: dataA <= 32'b00001111010000111011011001101000;
11'b01100100010: dataA <= 32'b10010110101000111101001101101001;
11'b01100100011: dataA <= 32'b00000001010101100000111010000001;
11'b01100100100: dataA <= 32'b01011000000100001100000011001110;
11'b01100100101: dataA <= 32'b00000001010000010100110000010010;
11'b01100100110: dataA <= 32'b01101100001010001000010100110001;
11'b01100100111: dataA <= 32'b00000110011010100011100000111010;
11'b01100101000: dataA <= 32'b10010100110001111011000110010000;
11'b01100101001: dataA <= 32'b00001001000100100000101101001001;
11'b01100101010: dataA <= 32'b11100011101100101110101100101111;
11'b01100101011: dataA <= 32'b00000110000001011000100010101101;
11'b01100101100: dataA <= 32'b01110010111100100110011000110001;
11'b01100101101: dataA <= 32'b00000000110000100010011010001101;
11'b01100101110: dataA <= 32'b10101100101010101101111111010001;
11'b01100101111: dataA <= 32'b00000101001001011110011110001011;
11'b01100110000: dataA <= 32'b00010010111000001100100100010001;
11'b01100110001: dataA <= 32'b00000100010010100110110100011011;
11'b01100110010: dataA <= 32'b10010101000010011001010010010001;
11'b01100110011: dataA <= 32'b00000110011011110101100010011001;
11'b01100110100: dataA <= 32'b11100101111000111111000111011001;
11'b01100110101: dataA <= 32'b00000011010011101110100110100100;
11'b01100110110: dataA <= 32'b10011000110110100011001101101010;
11'b01100110111: dataA <= 32'b00001010101111110110111101000010;
11'b01100111000: dataA <= 32'b00010110101011001101000111111110;
11'b01100111001: dataA <= 32'b00000011101101100100010100110011;
11'b01100111010: dataA <= 32'b01011100010000110100100101110000;
11'b01100111011: dataA <= 32'b00000110111000101111001000101001;
11'b01100111100: dataA <= 32'b01101101100111011100001111010011;
11'b01100111101: dataA <= 32'b00000001101011011110101011001101;
11'b01100111110: dataA <= 32'b10010101011101100111101011110111;
11'b01100111111: dataA <= 32'b00000110001110100010110011011010;
11'b01101000000: dataA <= 32'b01011110100101010110001110001110;
11'b01101000001: dataA <= 32'b00000111010110011101111000011100;
11'b01101000010: dataA <= 32'b00100111011010011100011100001110;
11'b01101000011: dataA <= 32'b00001111001111111101000101101110;
11'b01101000100: dataA <= 32'b00010111000101100111001000111110;
11'b01101000101: dataA <= 32'b00001010000001011110111111000001;
11'b01101000110: dataA <= 32'b11110000101110001101101011110101;
11'b01101000111: dataA <= 32'b00001110010001101101101100011101;
11'b01101001000: dataA <= 32'b11111001001111000100001110110010;
11'b01101001001: dataA <= 32'b00000011101100100100100111110011;
11'b01101001010: dataA <= 32'b00011011110001110010111100000101;
11'b01101001011: dataA <= 32'b00001010101000011011000101111101;
11'b01101001100: dataA <= 32'b10111100111000001011011011000010;
11'b01101001101: dataA <= 32'b00000100010001011010111110111100;
11'b01101001110: dataA <= 32'b11110110100101010101111100101101;
11'b01101001111: dataA <= 32'b00000111010100101110111001100100;
11'b01101010000: dataA <= 32'b10011110110010100000011010000110;
11'b01101010001: dataA <= 32'b00000010000110010100011000001100;
11'b01101010010: dataA <= 32'b01100011111010011101111101010100;
11'b01101010011: dataA <= 32'b00001111010001011001111010101110;
11'b01101010100: dataA <= 32'b01111001011110101100110111011011;
11'b01101010101: dataA <= 32'b00000001101110101000011010110101;
11'b01101010110: dataA <= 32'b00011100110101110000010110000101;
11'b01101010111: dataA <= 32'b00000011110101011011001101010100;
11'b01101011000: dataA <= 32'b10011110011101111001010010001110;
11'b01101011001: dataA <= 32'b00000111011101100101101010111000;
11'b01101011010: dataA <= 32'b00000000000011001010011010101101;
11'b01101011011: dataA <= 32'b00000000000000000000000000000000;
11'b01101011100: dataA <= 32'b11101010010001100000011001000001;
11'b01101011101: dataA <= 32'b00000101110100100110100100110110;
11'b01101011110: dataA <= 32'b00111101000000001100010010101101;
11'b01101011111: dataA <= 32'b00000111111110101011101111011011;
11'b01101100000: dataA <= 32'b10001110001110011110001011110101;
11'b01101100001: dataA <= 32'b00000100111101011111011000100001;
11'b01101100010: dataA <= 32'b00100010100001001001110110101010;
11'b01101100011: dataA <= 32'b00001011010001110100111000011110;
11'b01101100100: dataA <= 32'b00111010101001110101111001010011;
11'b01101100101: dataA <= 32'b00000111000110100110000101110111;
11'b01101100110: dataA <= 32'b01011100111000100110010100010011;
11'b01101100111: dataA <= 32'b00000110110110110110011001010100;
11'b01101101000: dataA <= 32'b11100111000010101101101101110101;
11'b01101101001: dataA <= 32'b00001100001010011111101001111100;
11'b01101101010: dataA <= 32'b00000111000011001101101111010010;
11'b01101101011: dataA <= 32'b00000110011110101101000000011010;
11'b01101101100: dataA <= 32'b00001111001100101100100101110000;
11'b01101101101: dataA <= 32'b00001011100011011001011001011001;
11'b01101101110: dataA <= 32'b00110011100110010111101111010001;
11'b01101101111: dataA <= 32'b00000111111000011011111010100111;
11'b01101110000: dataA <= 32'b01100110011010011110001100111011;
11'b01101110001: dataA <= 32'b00001000010110110010111010000000;
11'b01101110010: dataA <= 32'b10011010101010000011110110110101;
11'b01101110011: dataA <= 32'b00000101111110110100011101010011;
11'b01101110100: dataA <= 32'b11111010100100001100100001110111;
11'b01101110101: dataA <= 32'b00001000010100011101100110010101;
11'b01101110110: dataA <= 32'b11011100010110100011000111010111;
11'b01101110111: dataA <= 32'b00001111001010111101000101000000;
11'b01101111000: dataA <= 32'b10010010110001010101101100000101;
11'b01101111001: dataA <= 32'b00000010111010011110111001100001;
11'b01101111010: dataA <= 32'b11001100010000010101010011010001;
11'b01101111011: dataA <= 32'b00000010010101010010111100001011;
11'b01101111100: dataA <= 32'b00100000000101100000010101110011;
11'b01101111101: dataA <= 32'b00001000011011101001011100110011;
11'b01101111110: dataA <= 32'b01010010111101110011000110010001;
11'b01101111111: dataA <= 32'b00000110100100011110101100110010;
11'b01110000000: dataA <= 32'b01101011100101010111011100001100;
11'b01110000001: dataA <= 32'b00000011100011010010101010111101;
11'b01110000010: dataA <= 32'b00110000110001001111011000110001;
11'b01110000011: dataA <= 32'b00000001010101011010011110011101;
11'b01110000100: dataA <= 32'b01100110100010111101011110101011;
11'b01110000101: dataA <= 32'b00000011101011011000100010000011;
11'b01110000110: dataA <= 32'b01010011000100011101110100110100;
11'b01110000111: dataA <= 32'b00000100110101100100110000011100;
11'b01110001000: dataA <= 32'b10010101001001111001000010110110;
11'b01110001001: dataA <= 32'b00001000111011111011001101111001;
11'b01110001010: dataA <= 32'b01101111110001100111101001011000;
11'b01110001011: dataA <= 32'b00000011110110101000011110101100;
11'b01110001100: dataA <= 32'b01011000111010011010111100000110;
11'b01110001101: dataA <= 32'b00001010101101110100101100110011;
11'b01110001110: dataA <= 32'b00010010110011010100001010111101;
11'b01110001111: dataA <= 32'b00000011010001011100010100110100;
11'b01110010000: dataA <= 32'b10010100011001000101010110010010;
11'b01110010001: dataA <= 32'b00001000111001101110111100010010;
11'b01110010010: dataA <= 32'b01110011011011010011001111001110;
11'b01110010011: dataA <= 32'b00000001010000011010101011011100;
11'b01110010100: dataA <= 32'b10011011100110010111101100110011;
11'b01110010101: dataA <= 32'b00000110001111100000110011000001;
11'b01110010110: dataA <= 32'b01011000101001110110011101101010;
11'b01110010111: dataA <= 32'b00001000110110101001111000100101;
11'b01110011000: dataA <= 32'b01101011010010011100001011101011;
11'b01110011001: dataA <= 32'b00001110101001111100110010001110;
11'b01110011010: dataA <= 32'b10011001001110001111001011011101;
11'b01110011011: dataA <= 32'b00000111100001011110111110011000;
11'b01110011100: dataA <= 32'b11101100100010011101001100110010;
11'b01110011101: dataA <= 32'b00001110001100110101100000110110;
11'b01110011110: dataA <= 32'b01111000111011000011001110101101;
11'b01110011111: dataA <= 32'b00000011001111100000100011101010;
11'b01110100000: dataA <= 32'b00100101110001100011001001100010;
11'b01110100001: dataA <= 32'b00001001000110011101001010001101;
11'b01110100010: dataA <= 32'b11111010100000001100101000000001;
11'b01110100011: dataA <= 32'b00000100110100011011000010111011;
11'b01110100100: dataA <= 32'b00110000010101101110011011101010;
11'b01110100101: dataA <= 32'b00001000010100101100101101110101;
11'b01110100110: dataA <= 32'b11011100110101110000011000000101;
11'b01110100111: dataA <= 32'b00000000101011001110100100011101;
11'b01110101000: dataA <= 32'b10101101110110110101011101110000;
11'b01110101001: dataA <= 32'b00001111001011100011111011000101;
11'b01110101010: dataA <= 32'b10111101001010110100001001111011;
11'b01110101011: dataA <= 32'b00000001110011100000010110111100;
11'b01110101100: dataA <= 32'b10011010111001000000100100000111;
11'b01110101101: dataA <= 32'b00000101011000011101001101010100;
11'b01110101110: dataA <= 32'b01011000100001011001100010010011;
11'b01110101111: dataA <= 32'b00001001111101101101100010001000;
11'b01110110000: dataA <= 32'b00000000000010110001101010001011;
11'b01110110001: dataA <= 32'b00000000000000000000000000000000;
11'b01110110010: dataA <= 32'b10100000001000110001000110000001;
11'b01110110011: dataA <= 32'b00000110110101100000100001011111;
11'b01110110100: dataA <= 32'b00111100101000011101100010110001;
11'b01110110101: dataA <= 32'b00001010111110110011100111001010;
11'b01110110110: dataA <= 32'b00000110011110101101101100010001;
11'b01110110111: dataA <= 32'b00000111111110100011011000001011;
11'b01110111000: dataA <= 32'b00011100100000110010110101101100;
11'b01110111001: dataA <= 32'b00001011001111110010101000111111;
11'b01110111010: dataA <= 32'b11110100010110001101111001110010;
11'b01110111011: dataA <= 32'b00000101100111011100000110011110;
11'b01110111100: dataA <= 32'b11011100111001001111010101010110;
11'b01110111101: dataA <= 32'b00001000010111101100001001011100;
11'b01110111110: dataA <= 32'b11100110111010111100111110110000;
11'b01110111111: dataA <= 32'b00001010100111101001100110001100;
11'b01111000000: dataA <= 32'b10001001010011010100101110101100;
11'b01111000001: dataA <= 32'b00001001011110101100111000001011;
11'b01111000010: dataA <= 32'b11010011010100111101100110010010;
11'b01111000011: dataA <= 32'b00001000100001011111011100111001;
11'b01111000100: dataA <= 32'b01111001010111000111001111001011;
11'b01111000101: dataA <= 32'b00001001010111100111111011001110;
11'b01111000110: dataA <= 32'b01011110010110101101101110110111;
11'b01111000111: dataA <= 32'b00001001010101110000101001010000;
11'b01111001000: dataA <= 32'b00010110110010000011110111110110;
11'b01111001001: dataA <= 32'b00001000011110101100010001010100;
11'b01111001010: dataA <= 32'b10110010010000011110000011111100;
11'b01111001011: dataA <= 32'b00001001010100100101100110100101;
11'b01111001100: dataA <= 32'b11010100011010011010101000110111;
11'b01111001101: dataA <= 32'b00001101100101111100101100011001;
11'b01111001110: dataA <= 32'b00010000111101101110001001100011;
11'b01111001111: dataA <= 32'b00000101011101011110111001001010;
11'b01111010000: dataA <= 32'b01000100100000101110100011110101;
11'b01111010001: dataA <= 32'b00000011011001010011000100001101;
11'b01111010010: dataA <= 32'b00010100000100110001000110010101;
11'b01111010011: dataA <= 32'b00001010111010101111010100101100;
11'b01111010100: dataA <= 32'b01010011000101101011010110110010;
11'b01111010101: dataA <= 32'b00000100100110011010110000101011;
11'b01111010110: dataA <= 32'b01110001011010000111101011001001;
11'b01111010111: dataA <= 32'b00000001100111010000110111000100;
11'b01111011000: dataA <= 32'b10101100100101111111101000110000;
11'b01111011001: dataA <= 32'b00000010111010010100100010100100;
11'b01111011010: dataA <= 32'b01100000011111000100011101000110;
11'b01111011011: dataA <= 32'b00000011001111010010101001111011;
11'b01111011100: dataA <= 32'b01010101001100111111000101110110;
11'b01111011101: dataA <= 32'b00000110010111100000110000100101;
11'b01111011110: dataA <= 32'b10011001010001010001010100011001;
11'b01111011111: dataA <= 32'b00001011011010111010111001011001;
11'b01111100000: dataA <= 32'b11110111100010010111101010110111;
11'b01111100001: dataA <= 32'b00000101111001100000010110101011;
11'b01111100010: dataA <= 32'b01010111000010001010101010000011;
11'b01111100011: dataA <= 32'b00001001101011101110011100110100;
11'b01111100100: dataA <= 32'b00010000111111001011001101011010;
11'b01111100101: dataA <= 32'b00000011110100010100011000110101;
11'b01111100110: dataA <= 32'b00001110100101011110000110110011;
11'b01111100111: dataA <= 32'b00001010011000101100110000001100;
11'b01111101000: dataA <= 32'b01110101001011000010001110101000;
11'b01111101001: dataA <= 32'b00000001110101010110110011010011;
11'b01111101010: dataA <= 32'b11100011100110111111001101001111;
11'b01111101011: dataA <= 32'b00000110010001011100110010100000;
11'b01111101100: dataA <= 32'b01010100101110010110011100000110;
11'b01111101101: dataA <= 32'b00001001110101110011101100111110;
11'b01111101110: dataA <= 32'b00101101001010011011101010101000;
11'b01111101111: dataA <= 32'b00001101000101110110011010100110;
11'b01111110000: dataA <= 32'b10011101010010101110111101111001;
11'b01111110001: dataA <= 32'b00000100100010011110111101101000;
11'b01111110010: dataA <= 32'b10100100011010101100111100101110;
11'b01111110011: dataA <= 32'b00001100100111111001001101100111;
11'b01111110100: dataA <= 32'b01110110101010110010101101101000;
11'b01111110101: dataA <= 32'b00000011110011011010100111010001;
11'b01111110110: dataA <= 32'b11101111101001011011100111000010;
11'b01111110111: dataA <= 32'b00000111000110011111001010011100;
11'b01111111000: dataA <= 32'b00110010010000011110000101000001;
11'b01111111001: dataA <= 32'b00000101110110011011000110110011;
11'b01111111010: dataA <= 32'b01100110001110001110011010000111;
11'b01111111011: dataA <= 32'b00001001010100101000100110000101;
11'b01111111100: dataA <= 32'b00011010111001000000100101100110;
11'b01111111101: dataA <= 32'b00000000110000001010110000111111;
11'b01111111110: dataA <= 32'b11110111100110111100101101001100;
11'b01111111111: dataA <= 32'b00001101100110101111110111010100;
11'b10000000000: dataA <= 32'b11111010110010110011101011111001;
11'b10000000001: dataA <= 32'b00000011011000011000011011000011;
11'b10000000010: dataA <= 32'b00011010111100100001100010101010;
11'b10000000011: dataA <= 32'b00000111011001100001010001100101;
11'b10000000100: dataA <= 32'b01010010101001000010000011010111;
11'b10000000101: dataA <= 32'b00001100011010110011010101011000;
11'b10000000110: dataA <= 32'b00000000000010010001011001001010;
11'b10000000111: dataA <= 32'b00000000000000000000000000000000;
11'b10000001000: dataA <= 32'b00000100111100100110010000110011;
11'b10000001001: dataA <= 32'b00001010110010010000111111110101;
11'b10000001010: dataA <= 32'b10010100000110110111001000111010;
11'b10000001011: dataA <= 32'b00001111001010110010011001000001;
11'b10000001100: dataA <= 32'b10001111110010110010101000100111;
11'b10000001101: dataA <= 32'b00001111010000101100111001100111;
11'b10000001110: dataA <= 32'b00010001000101011110010110010100;
11'b10000001111: dataA <= 32'b00000111101001010100011011100110;
11'b10000010000: dataA <= 32'b00001010010110111011101001001100;
11'b10000010001: dataA <= 32'b00000011110100000011000111011011;
11'b10000010010: dataA <= 32'b00011101000111101101101011010101;
11'b10000010011: dataA <= 32'b00001011101111000100100110011101;
11'b10000010100: dataA <= 32'b10011100110010011010001000000010;
11'b10000010101: dataA <= 32'b00000011101010110010101110011011;
11'b10000010110: dataA <= 32'b10101001101110010001010110000010;
11'b10000010111: dataA <= 32'b00001111001101011100100101110111;
11'b10000011000: dataA <= 32'b00101011011010110110001001010011;
11'b10000011001: dataA <= 32'b00000000101110101111000000111110;
11'b10000011010: dataA <= 32'b10101010001111100001110101100001;
11'b10000011011: dataA <= 32'b00001011101101111100110011001001;
11'b10000011100: dataA <= 32'b01001011000010110010101011100010;
11'b10000011101: dataA <= 32'b00001010101101010100011100001101;
11'b10000011110: dataA <= 32'b01011001010001111011111011010000;
11'b10000011111: dataA <= 32'b00001111001111001000100110000101;
11'b10000100000: dataA <= 32'b11001000011011000111001110011000;
11'b10000100001: dataA <= 32'b00001010001101110010110110110010;
11'b10000100010: dataA <= 32'b00001101010101010011001011101110;
11'b10000100011: dataA <= 32'b00000010100100010110000100111111;
11'b10000100100: dataA <= 32'b10011111011111000100100001101100;
11'b10000100101: dataA <= 32'b00001110110101011101000001000101;
11'b10000100110: dataA <= 32'b10010001110111010110101010111000;
11'b10000100111: dataA <= 32'b00001100111001100011011010101111;
11'b10000101000: dataA <= 32'b10000011010100100110011010110011;
11'b10000101001: dataA <= 32'b00001101001010101010100010000110;
11'b10000101010: dataA <= 32'b10100011011001101100101001010010;
11'b10000101011: dataA <= 32'b00000011010110011001001001101110;
11'b10000101100: dataA <= 32'b11101100011111110011110100101001;
11'b10000101101: dataA <= 32'b00000011111100011011011110001001;
11'b10000101110: dataA <= 32'b11010010100111110100001000001110;
11'b10000101111: dataA <= 32'b00001101011010010001010110010010;
11'b10000110000: dataA <= 32'b00001110111110001001110011000101;
11'b10000110001: dataA <= 32'b00000111111001010101011001101100;
11'b10000110010: dataA <= 32'b11100111010111100110001011010100;
11'b10000110011: dataA <= 32'b00001011110011011000111110101110;
11'b10000110100: dataA <= 32'b00101001001100101101011100110111;
11'b10000110101: dataA <= 32'b00001101001001011100001000110101;
11'b10000110110: dataA <= 32'b10110000010011110011011011101010;
11'b10000110111: dataA <= 32'b00001100110100001010111101111010;
11'b10000111000: dataA <= 32'b01100001010001010011100001101011;
11'b10000111001: dataA <= 32'b00000101101100001110100010001110;
11'b10000111010: dataA <= 32'b01011111011101100001101101000101;
11'b10000111011: dataA <= 32'b00001010011000001101010110100110;
11'b10000111100: dataA <= 32'b10010011100011000101001001110010;
11'b10000111101: dataA <= 32'b00001100001011011000100110000111;
11'b10000111110: dataA <= 32'b01100100010101000001110100000010;
11'b10000111111: dataA <= 32'b00001010111100011001010001101001;
11'b10001000000: dataA <= 32'b11110010111011100010000111100101;
11'b10001000001: dataA <= 32'b00001000110011011001000100011010;
11'b10001000010: dataA <= 32'b00010111010111001011010011000111;
11'b10001000011: dataA <= 32'b00001010101100110110011011001110;
11'b10001000100: dataA <= 32'b11100100100101110011000100001010;
11'b10001000101: dataA <= 32'b00000010100101001100010011000010;
11'b10001000110: dataA <= 32'b10101001000111011010101100100100;
11'b10001000111: dataA <= 32'b00000001010110011111000000010100;
11'b10001001000: dataA <= 32'b11001100110110011010100111000110;
11'b10001001001: dataA <= 32'b00000011100110100110001111110100;
11'b10001001010: dataA <= 32'b01010100010001010010010100000100;
11'b10001001011: dataA <= 32'b00001001111000010011001000101001;
11'b10001001100: dataA <= 32'b00110100100001110101000001010001;
11'b10001001101: dataA <= 32'b00000011010001100101000010011011;
11'b10001001110: dataA <= 32'b01001000011011000111000000110101;
11'b10001001111: dataA <= 32'b00001011010100100011001001100010;
11'b10001010000: dataA <= 32'b11000110110011001011100011101011;
11'b10001010001: dataA <= 32'b00001010001101010010101110101011;
11'b10001010010: dataA <= 32'b00011101001000010101110011010100;
11'b10001010011: dataA <= 32'b00001000011110011001101011100110;
11'b10001010100: dataA <= 32'b01110010010010010010000110000101;
11'b10001010101: dataA <= 32'b00000011000100111010100010011001;
11'b10001010110: dataA <= 32'b11011000001001110010011100101000;
11'b10001010111: dataA <= 32'b00001100011001001101001101111001;
11'b10001011000: dataA <= 32'b11011111001000110110110101011010;
11'b10001011001: dataA <= 32'b00001100110001101000111110100100;
11'b10001011010: dataA <= 32'b00010101011001000101111011111001;
11'b10001011011: dataA <= 32'b00001101000111101010011000001101;
11'b10001011100: dataA <= 32'b00000000000000101011010101001101;
11'b10001011101: dataA <= 32'b00000000000000000000000000000000;
11'b10001011110: dataA <= 32'b01001000101000001100110000101101;
11'b10001011111: dataA <= 32'b00001010010100010010110011011110;
11'b10001100000: dataA <= 32'b00100000000110001111100110111010;
11'b10001100001: dataA <= 32'b00001111010000110110101001100001;
11'b10001100010: dataA <= 32'b11000111100011000011001010101000;
11'b10001100011: dataA <= 32'b00001110110110101101000000110110;
11'b10001100100: dataA <= 32'b00010000111000111101100101010010;
11'b10001100101: dataA <= 32'b00001000101001011100010111000111;
11'b10001100110: dataA <= 32'b01010100001010111100011001101101;
11'b10001100111: dataA <= 32'b00000011010001000010110011100100;
11'b10001101000: dataA <= 32'b01011101000111001110111001110111;
11'b10001101001: dataA <= 32'b00001011010010001100010010001101;
11'b10001101010: dataA <= 32'b00100000110010110010101010100100;
11'b10001101011: dataA <= 32'b00000101000111110101000010011100;
11'b10001101100: dataA <= 32'b00100001110010110001101001000001;
11'b10001101101: dataA <= 32'b00001111010011100000100101000111;
11'b10001101110: dataA <= 32'b00100111100010010110101000010100;
11'b10001101111: dataA <= 32'b00000001101000101101001100100101;
11'b10001110000: dataA <= 32'b11110010011011110011011000100001;
11'b10001110001: dataA <= 32'b00001100010000111101001011100010;
11'b10001110010: dataA <= 32'b11001100110011000011001101100110;
11'b10001110011: dataA <= 32'b00001011001111011100011000001011;
11'b10001110100: dataA <= 32'b01010101001001111011111010110010;
11'b10001110101: dataA <= 32'b00001111010100001110010101110101;
11'b10001110110: dataA <= 32'b01010010001010010111101011111100;
11'b10001110111: dataA <= 32'b00001010001111110011000110111011;
11'b10001111000: dataA <= 32'b11001011000101100010111011110001;
11'b10001111001: dataA <= 32'b00000101000001100010000100011101;
11'b10001111010: dataA <= 32'b11011001011010110101010010100111;
11'b10001111011: dataA <= 32'b00001101011010011101000000110100;
11'b10001111100: dataA <= 32'b10001001100110101111011000111001;
11'b10001111101: dataA <= 32'b00001010111011011111011001111111;
11'b10001111110: dataA <= 32'b01000010111100001100111001110100;
11'b10001111111: dataA <= 32'b00001101101111101110101101100110;
11'b10010000000: dataA <= 32'b01011111011001100100011000110011;
11'b10010000001: dataA <= 32'b00000010010010010111000001001110;
11'b10010000010: dataA <= 32'b00110010101011101101010110000111;
11'b10010000011: dataA <= 32'b00000001111000010101011010101010;
11'b10010000100: dataA <= 32'b00011000011111101101101000101110;
11'b10010000101: dataA <= 32'b00001010111101001111001010100011;
11'b10010000110: dataA <= 32'b11010000110010101010000101100010;
11'b10010000111: dataA <= 32'b00000101111000010001001101101011;
11'b10010001000: dataA <= 32'b00100011011010111111001010010110;
11'b10010001001: dataA <= 32'b00001010110110011000110110001111;
11'b10010001010: dataA <= 32'b00100101010100100100001011011010;
11'b10010001011: dataA <= 32'b00001101101110100110001000110100;
11'b10010001100: dataA <= 32'b10111000100011110100111100001101;
11'b10010001101: dataA <= 32'b00001011011000001110101110001010;
11'b10010001110: dataA <= 32'b01011101001101011011000011000111;
11'b10010001111: dataA <= 32'b00000110101010010110010101101110;
11'b10010010000: dataA <= 32'b01011001011010000001011110101010;
11'b10010010001: dataA <= 32'b00001000111001001011000110000110;
11'b10010010010: dataA <= 32'b01001101010110101101111001010011;
11'b10010010011: dataA <= 32'b00001100101110011110100001010111;
11'b10010010100: dataA <= 32'b00101100011001100001010111000001;
11'b10010010101: dataA <= 32'b00001000011101010101001010001001;
11'b10010010110: dataA <= 32'b11110011001011110011011001100110;
11'b10010010111: dataA <= 32'b00000111110011011000111100110001;
11'b10010011000: dataA <= 32'b11010101001111001100010101000100;
11'b10010011001: dataA <= 32'b00001011001110111100101110101110;
11'b10010011010: dataA <= 32'b10101000101010000011000101101000;
11'b10010011011: dataA <= 32'b00000100100010011000000111001011;
11'b10010011100: dataA <= 32'b00100111001111100011101110101001;
11'b10010011101: dataA <= 32'b00000000110000011111000000010011;
11'b10010011110: dataA <= 32'b01010000100110100011001001000110;
11'b10010011111: dataA <= 32'b00000110000011110000010111011110;
11'b10010100000: dataA <= 32'b10011100001101100001110110100010;
11'b10010100001: dataA <= 32'b00000111111001010000111101001000;
11'b10010100010: dataA <= 32'b10111000110101100100110001001100;
11'b10010100011: dataA <= 32'b00000011001101100101000110100011;
11'b10010100100: dataA <= 32'b00010000001010010111100000101111;
11'b10010100101: dataA <= 32'b00001010010110100001001001111010;
11'b10010100110: dataA <= 32'b01001010011111001100100101001000;
11'b10010100111: dataA <= 32'b00001010001111010110100110100100;
11'b10010101000: dataA <= 32'b00011011000100001100010010101111;
11'b10010101001: dataA <= 32'b00000101111110010011100010111111;
11'b10010101010: dataA <= 32'b11111010100110101010011000000100;
11'b10010101011: dataA <= 32'b00000101100001111100111010110001;
11'b10010101100: dataA <= 32'b00100100000110000010011101101100;
11'b10010101101: dataA <= 32'b00001001111100001010111110010010;
11'b10010101110: dataA <= 32'b01011101001000010101110011110111;
11'b10010101111: dataA <= 32'b00001100010101100111000110010101;
11'b10010110000: dataA <= 32'b10010001001100110101001001111011;
11'b10010110001: dataA <= 32'b00001110101100110000100100001011;
11'b10010110010: dataA <= 32'b00000000000000110010010101101011;
11'b10010110011: dataA <= 32'b00000000000000000000000000000000;
11'b10010110100: dataA <= 32'b01001110011000001011100001101000;
11'b10010110101: dataA <= 32'b00001001010101010110101010110111;
11'b10010110110: dataA <= 32'b00101100001001011111010100111000;
11'b10010110111: dataA <= 32'b00001110110110111010111110001001;
11'b10010111000: dataA <= 32'b11000011001111000100001011101010;
11'b10010111001: dataA <= 32'b00001100111011101011001100011101;
11'b10010111010: dataA <= 32'b10010010101100110100110101010000;
11'b10010111011: dataA <= 32'b00001001101011100100010110011111;
11'b10010111100: dataA <= 32'b01011110000110110101001010001111;
11'b10010111101: dataA <= 32'b00000011101101001000011011011101;
11'b10010111110: dataA <= 32'b01011011000010100111101000011000;
11'b10010111111: dataA <= 32'b00001010110100010110000101110101;
11'b10011000000: dataA <= 32'b01100010110010111011011100100111;
11'b10011000001: dataA <= 32'b00000111000110110011010010011100;
11'b10011000010: dataA <= 32'b01010111101111001010011011100011;
11'b10011000011: dataA <= 32'b00001110011000100110101000100110;
11'b10011000100: dataA <= 32'b11011111100001110110100111110100;
11'b10011000101: dataA <= 32'b00000011000100101001010100011011;
11'b10011000110: dataA <= 32'b00111000101111110100101011000010;
11'b10011000111: dataA <= 32'b00001011110011111001011111101100;
11'b10011001000: dataA <= 32'b01001110100111000100001111001100;
11'b10011001001: dataA <= 32'b00001011010001100010011000010010;
11'b10011001010: dataA <= 32'b00010101000001111011111010010100;
11'b10011001011: dataA <= 32'b00001101111001011000001001100101;
11'b10011001100: dataA <= 32'b00011100000101101111101001011110;
11'b10011001101: dataA <= 32'b00001010010001110001010110111100;
11'b10011001110: dataA <= 32'b10001010110101110010011011010100;
11'b10011001111: dataA <= 32'b00001000000001101100001000001100;
11'b10011010000: dataA <= 32'b11010101010010100110000100100100;
11'b10011010001: dataA <= 32'b00001010111101011100111100110011;
11'b10011010010: dataA <= 32'b01000011001110000111100111011001;
11'b10011010011: dataA <= 32'b00001000011101011001010101001111;
11'b10011010100: dataA <= 32'b00000100100100001011101000110110;
11'b10011010101: dataA <= 32'b00001101010011110000111001001110;
11'b10011010110: dataA <= 32'b10011001010101100100001000010011;
11'b10011010111: dataA <= 32'b00000010001101010110111100110101;
11'b10011011000: dataA <= 32'b10110110111011010110100111100110;
11'b10011011001: dataA <= 32'b00000000110011010001001110111010;
11'b10011011010: dataA <= 32'b10011110011011001110111000101110;
11'b10011011011: dataA <= 32'b00001000011110001100111010101011;
11'b10011011100: dataA <= 32'b10010100100110111010101000100001;
11'b10011011101: dataA <= 32'b00000100110101001111000001110011;
11'b10011011110: dataA <= 32'b00011101011010010111101000110111;
11'b10011011111: dataA <= 32'b00001001010111011010110001100111;
11'b10011100000: dataA <= 32'b00100001010100101011001000111011;
11'b10011100001: dataA <= 32'b00001101110011110000010100110011;
11'b10011100010: dataA <= 32'b11111100110111100110001100110001;
11'b10011100011: dataA <= 32'b00001001111001010010100010011010;
11'b10011100100: dataA <= 32'b11011011001101100010110101000100;
11'b10011100101: dataA <= 32'b00000111101010011110010001010101;
11'b10011100110: dataA <= 32'b01010101010010100001101111010000;
11'b10011100111: dataA <= 32'b00000110111000001010110101100110;
11'b10011101000: dataA <= 32'b10001001000110010110011000010100;
11'b10011101001: dataA <= 32'b00001100010010100100100000101110;
11'b10011101010: dataA <= 32'b10110010100110000001001001100001;
11'b10011101011: dataA <= 32'b00000101111100010101000010101001;
11'b10011101100: dataA <= 32'b00101111010111110100111011101000;
11'b10011101101: dataA <= 32'b00000111010011011000111001010001;
11'b10011101110: dataA <= 32'b00010011000011000101010111000011;
11'b10011101111: dataA <= 32'b00001011010001111101000110001111;
11'b10011110000: dataA <= 32'b10101100110010001011000111000111;
11'b10011110001: dataA <= 32'b00000111100001100010000111000100;
11'b10011110010: dataA <= 32'b11100011010011100100111111001110;
11'b10011110011: dataA <= 32'b00000000101011011111000000100001;
11'b10011110100: dataA <= 32'b00010110011110110011101010101000;
11'b10011110101: dataA <= 32'b00001000100011110110100110111111;
11'b10011110110: dataA <= 32'b01100110001110000001111001000010;
11'b10011110111: dataA <= 32'b00000110011000010010110101111000;
11'b10011111000: dataA <= 32'b00111001001001011100010010100111;
11'b10011111001: dataA <= 32'b00000100001010100011001010100100;
11'b10011111010: dataA <= 32'b00011100000101101111100001001001;
11'b10011111011: dataA <= 32'b00001000110111011111001010010010;
11'b10011111100: dataA <= 32'b11010010010010111101010110100110;
11'b10011111101: dataA <= 32'b00001010010001011100100010011100;
11'b10011111110: dataA <= 32'b10011001000000001010110011001011;
11'b10011111111: dataA <= 32'b00000011011011001101010110010111;
11'b10100000000: dataA <= 32'b10111100111010111011001010000101;
11'b10100000001: dataA <= 32'b00001000100001111101001111001010;
11'b10100000010: dataA <= 32'b01101110001110011010101101110001;
11'b10100000011: dataA <= 32'b00000111011100001100101110101010;
11'b10100000100: dataA <= 32'b01011011000100001100010010110011;
11'b10100000101: dataA <= 32'b00001010111000100111001010000101;
11'b10100000110: dataA <= 32'b00001111000000101100000111011011;
11'b10100000111: dataA <= 32'b00001110110001110100110100010010;
11'b10100001000: dataA <= 32'b00000000000001001001100110101010;
11'b10100001001: dataA <= 32'b00000000000000000000000000000000;
11'b10100001010: dataA <= 32'b10010110001100010010000011100011;
11'b10100001011: dataA <= 32'b00001000010110011010100110000111;
11'b10100001100: dataA <= 32'b01110100010100110110100011010101;
11'b10100001101: dataA <= 32'b00001101011011111001010010110001;
11'b10100001110: dataA <= 32'b01000010110110111100111100001110;
11'b10100001111: dataA <= 32'b00001010011110101001010100001100;
11'b10100010000: dataA <= 32'b10010110100100101011110101001110;
11'b10100010001: dataA <= 32'b00001010101100101100011101101111;
11'b10100010010: dataA <= 32'b01101010001010100101101010010001;
11'b10100010011: dataA <= 32'b00000100001010010000001011000110;
11'b10100010100: dataA <= 32'b00011010111101111111100110110111;
11'b10100010101: dataA <= 32'b00001001110110100000000101100101;
11'b10100010110: dataA <= 32'b10100100110111000100001110001011;
11'b10100010111: dataA <= 32'b00001001000110101111011110010100;
11'b10100011000: dataA <= 32'b11001111100011010011011101100111;
11'b10100011001: dataA <= 32'b00001100011100101010101100001100;
11'b10100011010: dataA <= 32'b11011001011101010110010110110011;
11'b10100011011: dataA <= 32'b00000110000001100101011000100010;
11'b10100011100: dataA <= 32'b01111011000011100110001101100110;
11'b10100011101: dataA <= 32'b00001010110110110001110011100101;
11'b10100011110: dataA <= 32'b01010110011010111100111111010001;
11'b10100011111: dataA <= 32'b00001010010100101010011100101001;
11'b10100100000: dataA <= 32'b10010100111001111011111001010101;
11'b10100100001: dataA <= 32'b00001011011101100010001001011100;
11'b10100100010: dataA <= 32'b11101000000100111111000110011110;
11'b10100100011: dataA <= 32'b00001001110011101011100010110100;
11'b10100100100: dataA <= 32'b00001110100110000010011010010110;
11'b10100100101: dataA <= 32'b00001011000010110110011000001011;
11'b10100100110: dataA <= 32'b11010011001010000110010111000011;
11'b10100100111: dataA <= 32'b00000111111110011100111100110010;
11'b10100101000: dataA <= 32'b10000010111001010111010101011000;
11'b10100101001: dataA <= 32'b00000101111100010101010000100110;
11'b10100101010: dataA <= 32'b00001010010000010010000111110110;
11'b10100101011: dataA <= 32'b00001100010111110001001000110101;
11'b10100101100: dataA <= 32'b10010101010001100011100111010011;
11'b10100101101: dataA <= 32'b00000011001001011000110100101100;
11'b10100101110: dataA <= 32'b10110101001010101111011001100111;
11'b10100101111: dataA <= 32'b00000000101101001111000011000011;
11'b10100110000: dataA <= 32'b00100110011110100111101000101111;
11'b10100110001: dataA <= 32'b00000101011101001110101110101100;
11'b10100110010: dataA <= 32'b10011010100011000011101011000011;
11'b10100110011: dataA <= 32'b00000011110010010000110101110011;
11'b10100110100: dataA <= 32'b01011001010101100111100111010111;
11'b10100110101: dataA <= 32'b00000111111000011110110000111110;
11'b10100110110: dataA <= 32'b01011101010100111010000110111011;
11'b10100110111: dataA <= 32'b00001100110111110110100101000010;
11'b10100111000: dataA <= 32'b01111011001111000111001100010100;
11'b10100111001: dataA <= 32'b00000111111010011010011010100011;
11'b10100111010: dataA <= 32'b00011001000101110010100111100010;
11'b10100111011: dataA <= 32'b00001000101010100110010100111101;
11'b10100111100: dataA <= 32'b11010011001010111010011110110101;
11'b10100111101: dataA <= 32'b00000101010111001110100101001101;
11'b10100111110: dataA <= 32'b01001010110101110110010111010100;
11'b10100111111: dataA <= 32'b00001011110101101000100100010101;
11'b10101000000: dataA <= 32'b01110100110110101001011100100100;
11'b10101000001: dataA <= 32'b00000011011001010100111011000010;
11'b10101000010: dataA <= 32'b10101001100011011110001100101100;
11'b10101000011: dataA <= 32'b00000110110010011010110101111000;
11'b10101000100: dataA <= 32'b11010010111010101110001001100100;
11'b10101000101: dataA <= 32'b00001010110011111011011101100110;
11'b10101000110: dataA <= 32'b01101110111110010011011001000111;
11'b10101000111: dataA <= 32'b00001010100001101110001010111101;
11'b10101001000: dataA <= 32'b00011111010111001110001111010100;
11'b10101001001: dataA <= 32'b00000010000110011111000001000001;
11'b10101001010: dataA <= 32'b10011110010110110100001100001011;
11'b10101001011: dataA <= 32'b00001010100100111000111010001111;
11'b10101001100: dataA <= 32'b01110000011010011010001011100100;
11'b10101001101: dataA <= 32'b00000100110110010100101010101000;
11'b10101001110: dataA <= 32'b10110101011101010011110100100100;
11'b10101001111: dataA <= 32'b00000101100111100001001010100100;
11'b10101010000: dataA <= 32'b01101000000100111111000010100101;
11'b10101010001: dataA <= 32'b00000111010111011101001010100010;
11'b10101010010: dataA <= 32'b00011100001110100110001000100110;
11'b10101010011: dataA <= 32'b00001001110011100010100010001101;
11'b10101010100: dataA <= 32'b10011000111100100001100100001000;
11'b10101010101: dataA <= 32'b00000001010110001011000101100111;
11'b10101010110: dataA <= 32'b10111101010011000011111100001000;
11'b10101010111: dataA <= 32'b00001011100010110111100111010011;
11'b10101011000: dataA <= 32'b00110110011110101010111101010110;
11'b10101011001: dataA <= 32'b00000101011011010010100010111011;
11'b10101011010: dataA <= 32'b01011011000000001010110010001111;
11'b10101011011: dataA <= 32'b00001000111001100011001101110101;
11'b10101011100: dataA <= 32'b00010000110100110010110100111010;
11'b10101011101: dataA <= 32'b00001101110110110101000100110001;
11'b10101011110: dataA <= 32'b00000000000001101001010111101001;
11'b10101011111: dataA <= 32'b00000000000000000000000000000000;
endcase
if (enB)
case(addrB)
11'b00000000000: dataB <= 32'b11000111010001000111010001111000;
11'b00000000001: dataB <= 32'b00001011001111010011001011110011;
11'b00000000010: dataB <= 32'b01001010010111010110011010111001;
11'b00000000011: dataB <= 32'b00001101100101101000001100101010;
11'b00000000100: dataB <= 32'b10011011111010011010000111000111;
11'b00000000101: dataB <= 32'b00001111001011101010101110001111;
11'b00000000110: dataB <= 32'b10010011010001111110100111010101;
11'b00000000111: dataB <= 32'b00000110001010001110100111110100;
11'b00000001000: dataB <= 32'b11000100101010110010111000101011;
11'b00000001001: dataB <= 32'b00000101010111000101011111001001;
11'b00000001010: dataB <= 32'b11011111001011110100001011110010;
11'b00000001011: dataB <= 32'b00001011001100000010111110100100;
11'b00000001100: dataB <= 32'b01011010110110000001110101100011;
11'b00000001101: dataB <= 32'b00000011001101101110100010010011;
11'b00000001110: dataB <= 32'b10110001100001101001010011100100;
11'b00000001111: dataB <= 32'b00001110000111010110101010011111;
11'b00000010000: dataB <= 32'b11101111001111001101011001110010;
11'b00000010001: dataB <= 32'b00000000110011101100110101011110;
11'b00000010010: dataB <= 32'b11100000001011000000110011000100;
11'b00000010011: dataB <= 32'b00001011001010111000011110101000;
11'b00000010100: dataB <= 32'b10001101010010011010001000100001;
11'b00000010101: dataB <= 32'b00001010001011001110101000101110;
11'b00000010110: dataB <= 32'b00011101010101111100001010101101;
11'b00000010111: dataB <= 32'b00001110101001000100111010010101;
11'b00000011000: dataB <= 32'b01000010101111100110001111010011;
11'b00000011001: dataB <= 32'b00001001101100110000101010011010;
11'b00000011010: dataB <= 32'b10010011100001001011111011001011;
11'b00000011011: dataB <= 32'b00000001001001001100010001100111;
11'b00000011100: dataB <= 32'b01100101011011001011110001110001;
11'b00000011101: dataB <= 32'b00001111010000011111000101011110;
11'b00000011110: dataB <= 32'b11011101111011101101011100010101;
11'b00000011111: dataB <= 32'b00001110010100101001010111010110;
11'b00000100000: dataB <= 32'b01001001101001000111011011010000;
11'b00000100001: dataB <= 32'b00001011100111100100011110100110;
11'b00000100010: dataB <= 32'b10101001010101110100111001110001;
11'b00000100011: dataB <= 32'b00000100111001011011001110010110;
11'b00000100100: dataB <= 32'b11100100010111101010100011101100;
11'b00000100101: dataB <= 32'b00000110111110100001100001110001;
11'b00000100110: dataB <= 32'b10001110110011110010110111101110;
11'b00000100111: dataB <= 32'b00001110110101010111100010000010;
11'b00000101000: dataB <= 32'b01010001001001110001110001101001;
11'b00000101001: dataB <= 32'b00001001011000011011011101110100;
11'b00000101010: dataB <= 32'b00101011001111110100111011110001;
11'b00000101011: dataB <= 32'b00001100010000011001000011001110;
11'b00000101100: dataB <= 32'b11101011000101000110001101110010;
11'b00000101101: dataB <= 32'b00001011100110010010010001001101;
11'b00000101110: dataB <= 32'b11100110001011100001111010000111;
11'b00000101111: dataB <= 32'b00001101010000001101001001101010;
11'b00000110000: dataB <= 32'b00100011001101010100010001010000;
11'b00000110001: dataB <= 32'b00000101001110001010110010100110;
11'b00000110010: dataB <= 32'b10100101011001001010001010100010;
11'b00000110011: dataB <= 32'b00001011110101010011100010111101;
11'b00000110100: dataB <= 32'b01011011101011001100011010010001;
11'b00000110101: dataB <= 32'b00001010101000010010101110101111;
11'b00000110110: dataB <= 32'b11011010010100101010100010000110;
11'b00000110111: dataB <= 32'b00001100111001011101010101001001;
11'b00000111000: dataB <= 32'b00110000101111000001000110000110;
11'b00000111001: dataB <= 32'b00001001010010011011001000010100;
11'b00000111010: dataB <= 32'b11011101011011000010100010001100;
11'b00000111011: dataB <= 32'b00001001101010101110001011011100;
11'b00000111100: dataB <= 32'b00011110100001101011010011101101;
11'b00000111101: dataB <= 32'b00000000101010000100100010101010;
11'b00000111110: dataB <= 32'b11101011000011000001101010000001;
11'b00000111111: dataB <= 32'b00000011011011100001000000100101;
11'b00001000000: dataB <= 32'b10001011000010000010010101100111;
11'b00001000001: dataB <= 32'b00000010001010011100001111110011;
11'b00001000010: dataB <= 32'b10001100011101000011000010001000;
11'b00001000011: dataB <= 32'b00001011010110010101010100001010;
11'b00001000100: dataB <= 32'b11101110010101111101010010010110;
11'b00001000101: dataB <= 32'b00000011110100100100111110010010;
11'b00001000110: dataB <= 32'b11000010101111100110000010111010;
11'b00001000111: dataB <= 32'b00001011110001100101000101001010;
11'b00001001000: dataB <= 32'b10000111000111000010110011001110;
11'b00001001001: dataB <= 32'b00001001101100010000111010100011;
11'b00001001010: dataB <= 32'b11011111001100110110110100010111;
11'b00001001011: dataB <= 32'b00001011011101100011101011110100;
11'b00001001100: dataB <= 32'b01101000000101111001110100000111;
11'b00001001101: dataB <= 32'b00000001001000110010010001110001;
11'b00001001110: dataB <= 32'b00001110010001011010101011000101;
11'b00001001111: dataB <= 32'b00001101110101010001011001100010;
11'b00001010000: dataB <= 32'b01100001001001011111100111111011;
11'b00001010001: dataB <= 32'b00001100101110100110111010101100;
11'b00001010010: dataB <= 32'b01011011011101011110011101010110;
11'b00001010011: dataB <= 32'b00001011000100100010010100100110;
11'b00001010100: dataB <= 32'b00000000000000101100100100110000;
11'b00001010101: dataB <= 32'b00000000000000000000000000000000;
11'b00001010110: dataB <= 32'b01001101100001110111100100011100;
11'b00001010111: dataB <= 32'b00001010101101010101010011101010;
11'b00001011000: dataB <= 32'b10000100100111101101001100010110;
11'b00001011001: dataB <= 32'b00001011000010011110001000100011;
11'b00001011010: dataB <= 32'b00100111111010000001110101001000;
11'b00001011011: dataB <= 32'b00001101100110100110101010111111;
11'b00001011100: dataB <= 32'b00010111011010011110011000010101;
11'b00001011101: dataB <= 32'b00000101101100001010110111110011;
11'b00001011110: dataB <= 32'b00000011000010100010010111101011;
11'b00001011111: dataB <= 32'b00000110111000001101101110101001;
11'b00001100000: dataB <= 32'b01100001001011110010111100001111;
11'b00001100001: dataB <= 32'b00001010001010000011010010101100;
11'b00001100010: dataB <= 32'b00011000111001101010000011100110;
11'b00001100011: dataB <= 32'b00000011010001101000011010001011;
11'b00001100100: dataB <= 32'b11110111010001001001100001101000;
11'b00001100101: dataB <= 32'b00001100000011010100110011001110;
11'b00001100110: dataB <= 32'b00110001000011010100011010010000;
11'b00001100111: dataB <= 32'b00000010011001101010101101111111;
11'b00001101000: dataB <= 32'b10010110001110010000010001001001;
11'b00001101001: dataB <= 32'b00001001101000101110001110000000;
11'b00001101010: dataB <= 32'b01010011100010000001110110000001;
11'b00001101011: dataB <= 32'b00001000101001001100111001001111;
11'b00001101100: dataB <= 32'b11100001010101111100001010001011;
11'b00001101101: dataB <= 32'b00001100100100000101001110100100;
11'b00001101110: dataB <= 32'b00000011000111110100101111001101;
11'b00001101111: dataB <= 32'b00001000101011101010011110000010;
11'b00001110000: dataB <= 32'b10011011101001001100011010001001;
11'b00001110001: dataB <= 32'b00000000101111000100100110010111;
11'b00001110010: dataB <= 32'b01101001010111000010110010010110;
11'b00001110011: dataB <= 32'b00001110101010011111000101111110;
11'b00001110100: dataB <= 32'b10100111111011110011111100110001;
11'b00001110101: dataB <= 32'b00001110101111101011001111101101;
11'b00001110110: dataB <= 32'b10010011110101110111101011001110;
11'b00001110111: dataB <= 32'b00001001100101011100011111000101;
11'b00001111000: dataB <= 32'b01101011001110000100111001101111;
11'b00001111001: dataB <= 32'b00000110111011011111010010110110;
11'b00001111010: dataB <= 32'b00011100010011010001010011010000;
11'b00001111011: dataB <= 32'b00001001111110100111011101010010;
11'b00001111100: dataB <= 32'b10001101000011011001100111001110;
11'b00001111101: dataB <= 32'b00001111001111011101100101110010;
11'b00001111110: dataB <= 32'b01010011010101010010000000101110;
11'b00001111111: dataB <= 32'b00001010110110100001100001110100;
11'b00010000000: dataB <= 32'b11101101000111110011011011101110;
11'b00010000001: dataB <= 32'b00001011101101011001001011100100;
11'b00010000010: dataB <= 32'b01101010111101100110101101101110;
11'b00010000011: dataB <= 32'b00001001100100001010011101100110;
11'b00010000100: dataB <= 32'b00011010000111000000111000100110;
11'b00010000101: dataB <= 32'b00001100101100010001011001011011;
11'b00010000110: dataB <= 32'b01100111001001011100110010010101;
11'b00010000111: dataB <= 32'b00000101010000001001000010111101;
11'b00010001000: dataB <= 32'b11101001010100110010111000000001;
11'b00010001001: dataB <= 32'b00001100010010011011101011001100;
11'b00010001010: dataB <= 32'b10100011101111001011011010001111;
11'b00010001011: dataB <= 32'b00001001000111010000110111010110;
11'b00010001100: dataB <= 32'b10010010011000100011110000101100;
11'b00010001101: dataB <= 32'b00001110010100100001010100110010;
11'b00010001110: dataB <= 32'b01101010100010011000010100001000;
11'b00010001111: dataB <= 32'b00001001110001011101001100100101;
11'b00010010000: dataB <= 32'b10100001011010101001110001110001;
11'b00010010001: dataB <= 32'b00001000101001100010000111100011;
11'b00010010010: dataB <= 32'b11011000100101100011100011110001;
11'b00010010011: dataB <= 32'b00000000110000000010111010010001;
11'b00010010100: dataB <= 32'b11101000111010011000110111000001;
11'b00010010101: dataB <= 32'b00000101111110100001000000111110;
11'b00010010110: dataB <= 32'b00001111010001110010010100001010;
11'b00010010111: dataB <= 32'b00000001101110010010010011100010;
11'b00010011000: dataB <= 32'b00000110110000111011110001001101;
11'b00010011001: dataB <= 32'b00001100010011011011011000001100;
11'b00010011010: dataB <= 32'b11100100001110001101000011111010;
11'b00010011011: dataB <= 32'b00000101010111100100111010000010;
11'b00010011100: dataB <= 32'b01000011000111110100100100111101;
11'b00010011101: dataB <= 32'b00001011101110100101000001000011;
11'b00010011110: dataB <= 32'b00001001011010101010000011010010;
11'b00010011111: dataB <= 32'b00001000101011010001000110011011;
11'b00010100000: dataB <= 32'b01100001001101011111100101111001;
11'b00010100001: dataB <= 32'b00001101111001101011100111110011;
11'b00010100010: dataB <= 32'b10011100000101100010000010101011;
11'b00010100011: dataB <= 32'b00000000101110100110000101010001;
11'b00010100100: dataB <= 32'b10000110100001010011001000100100;
11'b00010100101: dataB <= 32'b00001110010001010111100101001010;
11'b00010100110: dataB <= 32'b11100011001010001111101001111010;
11'b00010100111: dataB <= 32'b00001100001010100100110010101011;
11'b00010101000: dataB <= 32'b01100001100010000110101101110001;
11'b00010101001: dataB <= 32'b00001000100010011010010101000111;
11'b00010101010: dataB <= 32'b00000000000000110101100101010010;
11'b00010101011: dataB <= 32'b00000000000000000000000000000000;
11'b00010101100: dataB <= 32'b00010101101110011111100110111110;
11'b00010101101: dataB <= 32'b00001010001011011001011011001001;
11'b00010101110: dataB <= 32'b11000010111111110011101101010010;
11'b00010101111: dataB <= 32'b00001000000001010100010000100100;
11'b00010110000: dataB <= 32'b01110001110001100001110100001010;
11'b00010110001: dataB <= 32'b00001011000010100000100111011110;
11'b00010110010: dataB <= 32'b11011101011110110110001001010101;
11'b00010110011: dataB <= 32'b00000100101110001011000111100001;
11'b00010110100: dataB <= 32'b11000101010110001010000110101100;
11'b00010110101: dataB <= 32'b00001000111001011001111010001000;
11'b00010110110: dataB <= 32'b10100011000111011001101011101100;
11'b00010110111: dataB <= 32'b00001001001001001001100110101011;
11'b00010111000: dataB <= 32'b00011000111101010010010010001010;
11'b00010111001: dataB <= 32'b00000011110101100000010110000011;
11'b00010111010: dataB <= 32'b11111000111100110010010000101101;
11'b00010111011: dataB <= 32'b00001001100001010010111111100101;
11'b00010111100: dataB <= 32'b11110000110011010011011010001111;
11'b00010111101: dataB <= 32'b00000100011100100110100110100110;
11'b00010111110: dataB <= 32'b11001100011001101000010000101110;
11'b00010111111: dataB <= 32'b00001000000111100100000101011000;
11'b00011000000: dataB <= 32'b10011001100101100001110011000100;
11'b00011000001: dataB <= 32'b00000111101001001101000101111111;
11'b00011000010: dataB <= 32'b01100101010101111100001001001010;
11'b00011000011: dataB <= 32'b00001010000001001011100010101100;
11'b00011000100: dataB <= 32'b00000101011011110011011110001000;
11'b00011000101: dataB <= 32'b00000111101011100010011001101010;
11'b00011000110: dataB <= 32'b00100011101001011100111000101000;
11'b00011000111: dataB <= 32'b00000000110101000010111010111111;
11'b00011001000: dataB <= 32'b01101101001110101010010011111010;
11'b00011001001: dataB <= 32'b00001101000101100001000110011110;
11'b00011001010: dataB <= 32'b00110011101111101010101100101110;
11'b00011001011: dataB <= 32'b00001101101010101101000011110100;
11'b00011001100: dataB <= 32'b11011111111010011111101010001100;
11'b00011001101: dataB <= 32'b00000111100100010110100011001100;
11'b00011001110: dataB <= 32'b10101101000010001100111001101110;
11'b00011001111: dataB <= 32'b00001001011011100001010011001101;
11'b00011010000: dataB <= 32'b10010100011010101000100011110011;
11'b00011010001: dataB <= 32'b00001100011100101101010101000010;
11'b00011010010: dataB <= 32'b11001111001110110000100111001110;
11'b00011010011: dataB <= 32'b00001110101010100101100001100010;
11'b00011010100: dataB <= 32'b10011001011101000010100001010100;
11'b00011010101: dataB <= 32'b00001100010100100111011101111100;
11'b00011010110: dataB <= 32'b10101100111011100010001011001011;
11'b00011010111: dataB <= 32'b00001011001010011011001111100011;
11'b00011011000: dataB <= 32'b01101010110110000110111101001001;
11'b00011011001: dataB <= 32'b00000111000100000100110010000110;
11'b00011011010: dataB <= 32'b10010000001110011000010110100111;
11'b00011011011: dataB <= 32'b00001100001001010111100001010011;
11'b00011011100: dataB <= 32'b10100111000101100101000011111001;
11'b00011011101: dataB <= 32'b00000101010010001011010011001100;
11'b00011011110: dataB <= 32'b11101101001100101011110101000010;
11'b00011011111: dataB <= 32'b00001100101110100011101011001011;
11'b00011100000: dataB <= 32'b01101011100110111010101001101101;
11'b00011100001: dataB <= 32'b00000111000110010001000011101101;
11'b00011100010: dataB <= 32'b10001100100100101100110000110001;
11'b00011100011: dataB <= 32'b00001110101111100101010100100011;
11'b00011100100: dataB <= 32'b01100100011001101000010011001100;
11'b00011100101: dataB <= 32'b00001001110000011111001100111110;
11'b00011100110: dataB <= 32'b10100111010110001001100010010101;
11'b00011100111: dataB <= 32'b00000111001001010110000111011010;
11'b00011101000: dataB <= 32'b10010100101101100011110100010100;
11'b00011101001: dataB <= 32'b00000001010110000011001101110001;
11'b00011101010: dataB <= 32'b01100110110001110000110100100010;
11'b00011101011: dataB <= 32'b00001000011110100001000001100111;
11'b00011101100: dataB <= 32'b00010011011101100010110011001101;
11'b00011101101: dataB <= 32'b00000001110011001010011111001001;
11'b00011101110: dataB <= 32'b10000111000100111100110001010010;
11'b00011101111: dataB <= 32'b00001100110000011111011100010101;
11'b00011110000: dataB <= 32'b11011010001110011100110110011101;
11'b00011110001: dataB <= 32'b00000110111001100010110101110010;
11'b00011110010: dataB <= 32'b00000101011111110011010111111110;
11'b00011110011: dataB <= 32'b00001011001011100100111101000100;
11'b00011110100: dataB <= 32'b11001111101010010001100100010101;
11'b00011110101: dataB <= 32'b00000111101011010011010010001010;
11'b00011110110: dataB <= 32'b00100011001010001111100111111010;
11'b00011110111: dataB <= 32'b00001111010100110001011011100010;
11'b00011111000: dataB <= 32'b01010010001001001010100010001111;
11'b00011111001: dataB <= 32'b00000000110100011100000100111010;
11'b00011111010: dataB <= 32'b01000010110101001011110110000100;
11'b00011111011: dataB <= 32'b00001110001100011111101001000011;
11'b00011111100: dataB <= 32'b01100101000110111111011011111000;
11'b00011111101: dataB <= 32'b00001010100111100010110010101011;
11'b00011111110: dataB <= 32'b10100111011110100110011101101100;
11'b00011111111: dataB <= 32'b00000110000010010010011101110111;
11'b00100000000: dataB <= 32'b00000000000001001110010101110100;
11'b00100000001: dataB <= 32'b00000000000000000000000000000000;
11'b00100000010: dataB <= 32'b01011111110111001110111001111110;
11'b00100000011: dataB <= 32'b00001001001010011111011110100000;
11'b00100000100: dataB <= 32'b11000011010111100010011101001110;
11'b00100000101: dataB <= 32'b00000101000001001100011000110101;
11'b00100000110: dataB <= 32'b11111001100001010010010011101110;
11'b00100000111: dataB <= 32'b00001000000001011100100111110100;
11'b00100001000: dataB <= 32'b11100011011111001101001010010011;
11'b00100001001: dataB <= 32'b00000100110000001101010111000000;
11'b00100001010: dataB <= 32'b00001011101001110010000110001101;
11'b00100001011: dataB <= 32'b00001010011000100011111001100001;
11'b00100001100: dataB <= 32'b00100011000110110000101010101001;
11'b00100001101: dataB <= 32'b00000111101000010011110110100011;
11'b00100001110: dataB <= 32'b00011001000101000011000001001111;
11'b00100001111: dataB <= 32'b00000101011000010110011001110011;
11'b00100010000: dataB <= 32'b01110110101100101011010001010011;
11'b00100010001: dataB <= 32'b00000110100001010011000111110100;
11'b00100010010: dataB <= 32'b00101100101011000010011001101101;
11'b00100010011: dataB <= 32'b00000111011110100000100011000110;
11'b00100010100: dataB <= 32'b10000110101000111000110000110100;
11'b00100010101: dataB <= 32'b00000110101000011000000100110001;
11'b00100010110: dataB <= 32'b10100001101001010010010001001000;
11'b00100010111: dataB <= 32'b00000110101010001111010110101111;
11'b00100011000: dataB <= 32'b11101001001101111100001000001001;
11'b00100011001: dataB <= 32'b00000111100001010011101110101011;
11'b00100011010: dataB <= 32'b01001101101111100001111100000011;
11'b00100011011: dataB <= 32'b00000110101011011010011001011010;
11'b00100011100: dataB <= 32'b00101011100101100101010111001000;
11'b00100011101: dataB <= 32'b00000010011010000011010011100110;
11'b00100011110: dataB <= 32'b11101111000010010001110110011100;
11'b00100011111: dataB <= 32'b00001010100010100001000110110101;
11'b00100100000: dataB <= 32'b10111011011111010001011100001010;
11'b00100100001: dataB <= 32'b00001100100110101100111011110010;
11'b00100100010: dataB <= 32'b11101011111011001110111001101010;
11'b00100100011: dataB <= 32'b00000101000101010000101011010011;
11'b00100100100: dataB <= 32'b10101100111010010100101001001101;
11'b00100100101: dataB <= 32'b00001011011001100101001111010100;
11'b00100100110: dataB <= 32'b10001110100101111000010100110110;
11'b00100100111: dataB <= 32'b00001110011000101111001000111011;
11'b00100101000: dataB <= 32'b01010011011010000000010111001111;
11'b00100101001: dataB <= 32'b00001101000101101011011101011011;
11'b00100101010: dataB <= 32'b10011111100000111011100010111001;
11'b00100101011: dataB <= 32'b00001100110000101101010110000100;
11'b00100101100: dataB <= 32'b10101010110011000000111010001001;
11'b00100101101: dataB <= 32'b00001001101000011111001111011010;
11'b00100101110: dataB <= 32'b01100110101110101110101011100110;
11'b00100101111: dataB <= 32'b00000100100101000101000110100110;
11'b00100110000: dataB <= 32'b00001000011101101000010101001000;
11'b00100110001: dataB <= 32'b00001010000110011111101001010100;
11'b00100110010: dataB <= 32'b10101000111101110101010101111100;
11'b00100110011: dataB <= 32'b00000110010100010001100011001011;
11'b00100110100: dataB <= 32'b11101111000000110100110010100101;
11'b00100110101: dataB <= 32'b00001100001011101011100111001010;
11'b00100110110: dataB <= 32'b11110001011010100001111001001100;
11'b00100110111: dataB <= 32'b00000101100111010011001111110011;
11'b00100111000: dataB <= 32'b10001010110100111101110001010111;
11'b00100111001: dataB <= 32'b00001110001010101001001100101100;
11'b00100111010: dataB <= 32'b00011100011001000000110010110000;
11'b00100111011: dataB <= 32'b00001001101110100011001101011111;
11'b00100111100: dataB <= 32'b10101011010001101001100011111001;
11'b00100111101: dataB <= 32'b00000110001010001100010011000001;
11'b00100111110: dataB <= 32'b11010010110101100100010101010111;
11'b00100111111: dataB <= 32'b00000010111010001001100101011001;
11'b00101000000: dataB <= 32'b01100010101101010001000010000110;
11'b00101000001: dataB <= 32'b00001011011101100001000010010111;
11'b00101000010: dataB <= 32'b01011011100101010011000011010001;
11'b00101000011: dataB <= 32'b00000011011000000110110010011000;
11'b00101000100: dataB <= 32'b10001001010101001101010010010111;
11'b00101000101: dataB <= 32'b00001100001100100101011000101110;
11'b00101000110: dataB <= 32'b00010000010110100100011000111101;
11'b00101000111: dataB <= 32'b00001000111001100000110101100011;
11'b00101001000: dataB <= 32'b11001101101111100001111010111110;
11'b00101001001: dataB <= 32'b00001010001001100100111001001100;
11'b00101001010: dataB <= 32'b10011001110001110001100101111000;
11'b00101001011: dataB <= 32'b00000110101011010111011001111010;
11'b00101001100: dataB <= 32'b11100101000110111111011010011001;
11'b00101001101: dataB <= 32'b00001111001111110101001111000000;
11'b00101001110: dataB <= 32'b00001000011001000011010010110011;
11'b00101001111: dataB <= 32'b00000010011001010000001000101011;
11'b00101010000: dataB <= 32'b00000101001101001100010100000110;
11'b00101010001: dataB <= 32'b00001100100111100111100100111100;
11'b00101010010: dataB <= 32'b11100101000011011110011101010101;
11'b00101010011: dataB <= 32'b00001000100110011110101110011010;
11'b00101010100: dataB <= 32'b10101101010110111101111100101000;
11'b00101010101: dataB <= 32'b00000011100101001100101010100111;
11'b00101010110: dataB <= 32'b00000000000001101110100110110101;
11'b00101010111: dataB <= 32'b00000000000000000000000000000000;
11'b00101011000: dataB <= 32'b11111011000011011001101111001100;
11'b00101011001: dataB <= 32'b00000101001101101111000000001010;
11'b00101011010: dataB <= 32'b01101011111001001000110111000101;
11'b00101011011: dataB <= 32'b00000000110101001101100110111110;
11'b00101011100: dataB <= 32'b01110000001101001101010111011000;
11'b00101011101: dataB <= 32'b00000000101111010011000110011000;
11'b00101011110: dataB <= 32'b11101110111010100001101001101011;
11'b00101011111: dataB <= 32'b00001000010110101011100100011001;
11'b00101100000: dataB <= 32'b11110101101001000100010110110011;
11'b00101100001: dataB <= 32'b00001100001011111100111000100100;
11'b00101100010: dataB <= 32'b11100010111000010010010100101010;
11'b00101100011: dataB <= 32'b00000100010000111011011001100010;
11'b00101100100: dataB <= 32'b01100011001101100101110111111101;
11'b00101100101: dataB <= 32'b00001100010101001101010001100100;
11'b00101100110: dataB <= 32'b01010110010001101110101001111101;
11'b00101100111: dataB <= 32'b00000000110010100011011010001000;
11'b00101101000: dataB <= 32'b11010100100101001001110110101100;
11'b00101101001: dataB <= 32'b00001111010001010000111111000001;
11'b00101101010: dataB <= 32'b01010101110000011110001010011110;
11'b00101101011: dataB <= 32'b00000100010010000011001100110110;
11'b00101101100: dataB <= 32'b10110100111101001101010100011101;
11'b00101101101: dataB <= 32'b00000101010010101011100011110010;
11'b00101101110: dataB <= 32'b10100110101110000100000100101111;
11'b00101101111: dataB <= 32'b00000000110000110111011001111010;
11'b00101110000: dataB <= 32'b00110111100100111000110001100111;
11'b00101110001: dataB <= 32'b00000101110010001101001001001101;
11'b00101110010: dataB <= 32'b11110010101010101100110100010001;
11'b00101110011: dataB <= 32'b00001101011011101001111011000000;
11'b00101110100: dataB <= 32'b01100000100000111011011110010011;
11'b00101110101: dataB <= 32'b00000001001010100010111110111010;
11'b00101110110: dataB <= 32'b01101110001000101001010101000111;
11'b00101110111: dataB <= 32'b00000011000110011100100101010000;
11'b00101111000: dataB <= 32'b01111100101011011001100101001100;
11'b00101111001: dataB <= 32'b00000010110101010101011101111001;
11'b00101111010: dataB <= 32'b01011100100110010011010110101101;
11'b00101111011: dataB <= 32'b00001100101001100110110110010001;
11'b00101111100: dataB <= 32'b00010011100000001100001011010110;
11'b00101111101: dataB <= 32'b00001100000011100100100001110110;
11'b00101111110: dataB <= 32'b00101101011000001011110111110001;
11'b00101111111: dataB <= 32'b00000010100101101110101001101101;
11'b00110000000: dataB <= 32'b11110001000001110110001100111010;
11'b00110000001: dataB <= 32'b00001000000110101010100110010011;
11'b00110000010: dataB <= 32'b00011000101000011001110100101011;
11'b00110000011: dataB <= 32'b00000100001100100111000001010001;
11'b00110000100: dataB <= 32'b11010110110011010010100011001000;
11'b00110000101: dataB <= 32'b00000010110110100011110111001010;
11'b00110000110: dataB <= 32'b01001111101100001100100100010101;
11'b00110000111: dataB <= 32'b00000011001011110101000010000101;
11'b00110001000: dataB <= 32'b10011110101110101100011110010100;
11'b00110001001: dataB <= 32'b00001010010011110001011101110001;
11'b00110001010: dataB <= 32'b10100000100010011110010010111010;
11'b00110001011: dataB <= 32'b00000101100111110010101001011001;
11'b00110001100: dataB <= 32'b01101100011100111010110110001101;
11'b00110001101: dataB <= 32'b00000011110100100111011001111000;
11'b00110001110: dataB <= 32'b10011011101010111110001011111101;
11'b00110001111: dataB <= 32'b00000101000011100110101110010110;
11'b00110010000: dataB <= 32'b00001101000100011101111000011010;
11'b00110010001: dataB <= 32'b00000111001100100110111011100101;
11'b00110010010: dataB <= 32'b11101000101000110100101100111000;
11'b00110010011: dataB <= 32'b00000101010011001001100100110001;
11'b00110010100: dataB <= 32'b00011011011010001100111011110101;
11'b00110010101: dataB <= 32'b00001101011010110011101100111101;
11'b00110010110: dataB <= 32'b01010110111000100101010011011011;
11'b00110010111: dataB <= 32'b00001110101001100000111111101011;
11'b00110011000: dataB <= 32'b00110011001001100101011000111001;
11'b00110011001: dataB <= 32'b00001100011001011001110000001011;
11'b00110011010: dataB <= 32'b10101011101110101101101011111011;
11'b00110011011: dataB <= 32'b00000110000111101100110111010110;
11'b00110011100: dataB <= 32'b11001011011110001010111110101110;
11'b00110011101: dataB <= 32'b00001100101110011010111101100100;
11'b00110011110: dataB <= 32'b10110111100100111000111111001010;
11'b00110011111: dataB <= 32'b00000100101011011100110110011101;
11'b00110100000: dataB <= 32'b00111001001100110100011100010100;
11'b00110100001: dataB <= 32'b00000101110010101101010001010100;
11'b00110100010: dataB <= 32'b11100010110111101010001100101011;
11'b00110100011: dataB <= 32'b00000111100001100110010100011001;
11'b00110100100: dataB <= 32'b10001101101101101101111001111010;
11'b00110100101: dataB <= 32'b00001100111011000101011101100110;
11'b00110100110: dataB <= 32'b00100111110110001101100011010111;
11'b00110100111: dataB <= 32'b00000011100110110010110010000110;
11'b00110101000: dataB <= 32'b00100000110111001001001010100101;
11'b00110101001: dataB <= 32'b00000011001110010111000001011011;
11'b00110101010: dataB <= 32'b11101010100110111010000100000110;
11'b00110101011: dataB <= 32'b00000010111000010101100111110010;
11'b00110101100: dataB <= 32'b00000000000011010100101010110010;
11'b00110101101: dataB <= 32'b00000000000000000000000000000000;
11'b00110101110: dataB <= 32'b10110111010111110011001111010010;
11'b00110101111: dataB <= 32'b00000101101011101101001100100001;
11'b00110110000: dataB <= 32'b11011111111001110000011001000101;
11'b00110110001: dataB <= 32'b00000000101111001001010110011110;
11'b00110110010: dataB <= 32'b00111000011100111100110101010111;
11'b00110110011: dataB <= 32'b00000001001001010010111111001001;
11'b00110110100: dataB <= 32'b11101111000111000010011010101101;
11'b00110110101: dataB <= 32'b00000111010110100011101000111000;
11'b00110110110: dataB <= 32'b10101011110101000011100110010010;
11'b00110110111: dataB <= 32'b00001100101110111101001100011011;
11'b00110111000: dataB <= 32'b10100010111000110001000110001000;
11'b00110111001: dataB <= 32'b00000100101101110011101101110010;
11'b00110111010: dataB <= 32'b11011111001101001101010101011011;
11'b00110111011: dataB <= 32'b00001010111000001010111101100011;
11'b00110111100: dataB <= 32'b11011110001101001110010110111110;
11'b00110111101: dataB <= 32'b00000000101100011111011010111000;
11'b00110111110: dataB <= 32'b11011000011101101001010111101011;
11'b00110111111: dataB <= 32'b00001110010111010010110011011010;
11'b00111000000: dataB <= 32'b00001101100100001100100111011110;
11'b00111000001: dataB <= 32'b00000011101111000010110100011101;
11'b00111000010: dataB <= 32'b00110011001100111100110010011001;
11'b00111000011: dataB <= 32'b00000100110000100011100111110100;
11'b00111000100: dataB <= 32'b10101010110110000100000101001101;
11'b00111000101: dataB <= 32'b00000000101011110001101010001010;
11'b00111000110: dataB <= 32'b10101101110101101000010100000011;
11'b00111000111: dataB <= 32'b00000101110000001100111001000100;
11'b00111001000: dataB <= 32'b00110100111010011101000100001110;
11'b00111001001: dataB <= 32'b00001010111110011101111011100010;
11'b00111001010: dataB <= 32'b00100110100101001010101101011000;
11'b00111001011: dataB <= 32'b00000010100101100010111111001011;
11'b00111001100: dataB <= 32'b01110110011001010000100111000110;
11'b00111001101: dataB <= 32'b00000101000100100000100110000000;
11'b00111001110: dataB <= 32'b10111101000011110011000110001011;
11'b00111001111: dataB <= 32'b00000010010000010001010010011001;
11'b00111010000: dataB <= 32'b10100000100110011011100111001100;
11'b00111010001: dataB <= 32'b00001101101101101000111110110001;
11'b00111010010: dataB <= 32'b11001101010100010010101001111000;
11'b00111010011: dataB <= 32'b00001110000111101010100101010101;
11'b00111010100: dataB <= 32'b11100111100000010010010111010001;
11'b00111010101: dataB <= 32'b00000101000010110000110101011100;
11'b00111010110: dataB <= 32'b00101111001101010101111010011101;
11'b00111010111: dataB <= 32'b00001010000111101110110010010100;
11'b00111011000: dataB <= 32'b11011100100101000000110101101001;
11'b00111011001: dataB <= 32'b00000101001001100111001001110000;
11'b00111011010: dataB <= 32'b11011010101011011011110100100101;
11'b00111011011: dataB <= 32'b00000010010001011001110111001011;
11'b00111011100: dataB <= 32'b01000111011100001011000011110010;
11'b00111011101: dataB <= 32'b00000100100111110001010001110101;
11'b00111011110: dataB <= 32'b10100010110010100100111100111000;
11'b00111011111: dataB <= 32'b00001001010101101001101010010001;
11'b00111100000: dataB <= 32'b10100110100101111110100001010101;
11'b00111100001: dataB <= 32'b00000111000110110100111001111001;
11'b00111100010: dataB <= 32'b10110010101001010010000110101100;
11'b00111100011: dataB <= 32'b00000011010001100001011110101000;
11'b00111100100: dataB <= 32'b11010011100110011110101000111110;
11'b00111100101: dataB <= 32'b00000111100010101010110101110110;
11'b00111100110: dataB <= 32'b00001100110100001100100110011001;
11'b00111100111: dataB <= 32'b00001000001100100111000011001110;
11'b00111101000: dataB <= 32'b00101010110000110011101010111011;
11'b00111101001: dataB <= 32'b00000100110001000011010001010001;
11'b00111101010: dataB <= 32'b01010111010101111100111010010111;
11'b00111101011: dataB <= 32'b00001011011101100111111000110100;
11'b00111101100: dataB <= 32'b11011000110000011100010001010110;
11'b00111101101: dataB <= 32'b00001111001111100000111111101100;
11'b00111101110: dataB <= 32'b10101111011001011100110110111001;
11'b00111101111: dataB <= 32'b00001001111100001111101000100001;
11'b00111110000: dataB <= 32'b01100011110010011110001001011101;
11'b00111110001: dataB <= 32'b00001000000110101111000010110111;
11'b00111110010: dataB <= 32'b01000111001010011011001110110011;
11'b00111110011: dataB <= 32'b00001100110010011010111001011100;
11'b00111110100: dataB <= 32'b11101111110101101000011111010000;
11'b00111110101: dataB <= 32'b00000101101001011110110110000101;
11'b00111110110: dataB <= 32'b10110101100000110011011010110111;
11'b00111110111: dataB <= 32'b00000101110000101001011001011011;
11'b00111111000: dataB <= 32'b11100100111011110011101101010000;
11'b00111111001: dataB <= 32'b00001010000001101100011101000000;
11'b00111111010: dataB <= 32'b00000101011001010101100111111011;
11'b00111111011: dataB <= 32'b00001010011110000011000101001110;
11'b00111111100: dataB <= 32'b11011011111001111101100010010011;
11'b00111111101: dataB <= 32'b00000110000011110101000001101101;
11'b00111111110: dataB <= 32'b10100010110111101010001100001000;
11'b00111111111: dataB <= 32'b00000011101010011000111001101010;
11'b01000000000: dataB <= 32'b01101110110011001010110110000100;
11'b01000000001: dataB <= 32'b00000001010011001111011011110100;
11'b01000000010: dataB <= 32'b00000000000011001101101010010100;
11'b01000000011: dataB <= 32'b00000000000000000000000000000000;
11'b01000000100: dataB <= 32'b10110001100111110100011110010111;
11'b01000000101: dataB <= 32'b00000110101010101001010101001000;
11'b01000000110: dataB <= 32'b11010011110110100000101011000111;
11'b01000000111: dataB <= 32'b00000001001001000101000001110110;
11'b01000001000: dataB <= 32'b00111100110000111011110100010101;
11'b01000001001: dataB <= 32'b00000011000100010100110011100010;
11'b01000001010: dataB <= 32'b01101101010011001011001010101111;
11'b01000001011: dataB <= 32'b00000110010100011011101001100000;
11'b01000001100: dataB <= 32'b10100001111001001010110101110000;
11'b01000001101: dataB <= 32'b00001100010010110111100100100010;
11'b01000001110: dataB <= 32'b10100100111101011000010111100111;
11'b01000001111: dataB <= 32'b00000101001011101001111010001010;
11'b01000010000: dataB <= 32'b10011101001101000100100011011000;
11'b01000010001: dataB <= 32'b00001000111001001100101101100011;
11'b01000010010: dataB <= 32'b10101000010000110101100100011100;
11'b01000010011: dataB <= 32'b00000001100111011001010111011001;
11'b01000010100: dataB <= 32'b00100000011110001001011000001011;
11'b01000010101: dataB <= 32'b00001100111011010110101011100100;
11'b01000010110: dataB <= 32'b11000111010000001011010100111101;
11'b01000010111: dataB <= 32'b00000100001100000110100000010011;
11'b01000011000: dataB <= 32'b10110001011000111011110000110011;
11'b01000011001: dataB <= 32'b00000100101110011101100111101101;
11'b01000011010: dataB <= 32'b11101010111110000100000101101011;
11'b01000011011: dataB <= 32'b00000010000110100111110110011010;
11'b01000011100: dataB <= 32'b11100011111010010000010110100001;
11'b01000011101: dataB <= 32'b00000101101110001110101001000011;
11'b01000011110: dataB <= 32'b01110101001010001101100100101011;
11'b01000011111: dataB <= 32'b00000111111110010011110111110011;
11'b01000100000: dataB <= 32'b00101010101101011001111011011011;
11'b01000100001: dataB <= 32'b00000101000010100011000011001100;
11'b01000100010: dataB <= 32'b10111100110001111000011000100110;
11'b01000100011: dataB <= 32'b00000111100010100110101010110000;
11'b01000100100: dataB <= 32'b11111011011011110100010111001001;
11'b01000100101: dataB <= 32'b00000010101100001111000110110001;
11'b01000100110: dataB <= 32'b01100110101010011011110111101100;
11'b01000100111: dataB <= 32'b00001101110010101001000011001010;
11'b01000101000: dataB <= 32'b01001001000100101001011000011001;
11'b01000101001: dataB <= 32'b00001111001100101110110001000101;
11'b01000101010: dataB <= 32'b01100001100100110001000111010001;
11'b01000101011: dataB <= 32'b00000111100001110011000101010100;
11'b01000101100: dataB <= 32'b01101011011001000101010111011110;
11'b01000101101: dataB <= 32'b00001011001010110000111110001100;
11'b01000101110: dataB <= 32'b11100010100101101000010111001000;
11'b01000101111: dataB <= 32'b00000110101000100101001110011000;
11'b01000110000: dataB <= 32'b11011110101011010100110111000100;
11'b01000110001: dataB <= 32'b00000010001100001111101011001100;
11'b01000110010: dataB <= 32'b00000011001000011001110011001110;
11'b01000110011: dataB <= 32'b00000110000110101101011101100101;
11'b01000110100: dataB <= 32'b00100100110010011101001010111011;
11'b01000110101: dataB <= 32'b00001000010101100001101110101010;
11'b01000110110: dataB <= 32'b10101010101101011110010000101111;
11'b01000110111: dataB <= 32'b00001001000111110101001010011001;
11'b01000111000: dataB <= 32'b01110110111001101001100111101011;
11'b01000111001: dataB <= 32'b00000011101101011011011111010001;
11'b01000111010: dataB <= 32'b01001101011001111110110110011110;
11'b01000111011: dataB <= 32'b00001010000011101010111101010110;
11'b01000111100: dataB <= 32'b11010000101000001011000100010111;
11'b01000111101: dataB <= 32'b00001000101100100111000110101110;
11'b01000111110: dataB <= 32'b11101100111100111010101000111100;
11'b01000111111: dataB <= 32'b00000100101110000010111001110000;
11'b01001000000: dataB <= 32'b01010011001101110100111000111000;
11'b01001000001: dataB <= 32'b00001000011110011101111000111011;
11'b01001000010: dataB <= 32'b00011100101100011011000000110001;
11'b01001000011: dataB <= 32'b00001111010100100000111111011110;
11'b01001000100: dataB <= 32'b11101001100001001100010101010111;
11'b01001000101: dataB <= 32'b00000111011100001001011001000000;
11'b01001000110: dataB <= 32'b10011001110001111110000110111101;
11'b01001000111: dataB <= 32'b00001001100111101101001010000111;
11'b01001001000: dataB <= 32'b11000110110110100011101101011000;
11'b01001001001: dataB <= 32'b00001011110101011100110101011011;
11'b01001001010: dataB <= 32'b11100011111010010000011110110110;
11'b01001001011: dataB <= 32'b00000111001000100000110101101101;
11'b01001001100: dataB <= 32'b00101101101101000010101001011001;
11'b01001001101: dataB <= 32'b00000101101110100011011101100011;
11'b01001001110: dataB <= 32'b01100110111111110101001100110100;
11'b01001001111: dataB <= 32'b00001100100100110010101001101000;
11'b01001010000: dataB <= 32'b01000011000101000100110101111010;
11'b01001010001: dataB <= 32'b00000111011110000010110000110101;
11'b01001010010: dataB <= 32'b10010001110001100101010010001110;
11'b01001010011: dataB <= 32'b00001000100011110011010001010101;
11'b01001010100: dataB <= 32'b10100100111011110011101101001100;
11'b01001010101: dataB <= 32'b00000101000111011000110101111010;
11'b01001010110: dataB <= 32'b11110000111111010011111000100100;
11'b01001010111: dataB <= 32'b00000001001110001011001011101101;
11'b01001011000: dataB <= 32'b00000000000010110110011001010101;
11'b01001011001: dataB <= 32'b00000000000000000000000000000000;
11'b01001011010: dataB <= 32'b01101001110011101101111100011100;
11'b01001011011: dataB <= 32'b00000111101001100101011001111000;
11'b01001011100: dataB <= 32'b10001011101011001001011100101010;
11'b01001011101: dataB <= 32'b00000010100100000110101101001110;
11'b01001011110: dataB <= 32'b10111101001001000011000011110001;
11'b01001011111: dataB <= 32'b00000101100001010110101011110011;
11'b01001100000: dataB <= 32'b01101001011011010100001010110001;
11'b01001100001: dataB <= 32'b00000101010011010011100010010000;
11'b01001100010: dataB <= 32'b10010101110101011010010101101110;
11'b01001100011: dataB <= 32'b00001011110101101111110100111001;
11'b01001100100: dataB <= 32'b11100101000010000000011001001000;
11'b01001100101: dataB <= 32'b00000110001001011111111010011010;
11'b01001100110: dataB <= 32'b01011011001000111011110001110100;
11'b01001100111: dataB <= 32'b00000110111001010000100001101011;
11'b01001101000: dataB <= 32'b00110000011100101100100010011000;
11'b01001101001: dataB <= 32'b00000011100011010101010011110011;
11'b01001101010: dataB <= 32'b00100110100010101001101001001100;
11'b01001101011: dataB <= 32'b00001001111110011010100111011101;
11'b01001101100: dataB <= 32'b10000100111100011001110010011001;
11'b01001101101: dataB <= 32'b00000101001001001110001100011010;
11'b01001101110: dataB <= 32'b10101001100101000011000000101110;
11'b01001101111: dataB <= 32'b00000101101011010101100011010110;
11'b01001110000: dataB <= 32'b01101011000110000100000110101010;
11'b01001110001: dataB <= 32'b00000100100010011101110110100011;
11'b01001110010: dataB <= 32'b00010111111011000000111001100001;
11'b01001110011: dataB <= 32'b00000110001100010100011101001011;
11'b01001110100: dataB <= 32'b11110001011001111101100101101001;
11'b01001110101: dataB <= 32'b00000100111101001001100111110100;
11'b01001110110: dataB <= 32'b00101100110101111001101000111100;
11'b01001110111: dataB <= 32'b00001000000001100011000011001101;
11'b01001111000: dataB <= 32'b01111101000110101000101010100111;
11'b01001111001: dataB <= 32'b00001010000011101010101111011001;
11'b01001111010: dataB <= 32'b11110101101111101101111000001001;
11'b01001111011: dataB <= 32'b00000011101000001110110111001010;
11'b01001111100: dataB <= 32'b01101010101110011100011000101100;
11'b01001111101: dataB <= 32'b00001100110110100111001011010011;
11'b01001111110: dataB <= 32'b01001010110101010000100110011000;
11'b01001111111: dataB <= 32'b00001111010010110000111100111100;
11'b01010000000: dataB <= 32'b11011001100001011000010111010000;
11'b01010000001: dataB <= 32'b00001010100010110001010001010011;
11'b01010000010: dataB <= 32'b01100101011100111100010100111100;
11'b01010000011: dataB <= 32'b00001100001101101111001010001100;
11'b01010000100: dataB <= 32'b10100110101010011000011000101000;
11'b01010000101: dataB <= 32'b00001000000111100001001111000001;
11'b01010000110: dataB <= 32'b10100010101011000101111001000100;
11'b01010000111: dataB <= 32'b00000011001000001001011010111101;
11'b01010001000: dataB <= 32'b10000100110000111000110011101011;
11'b01010001001: dataB <= 32'b00001000000101100101100101011100;
11'b01010001010: dataB <= 32'b11100110111010001101011000011101;
11'b01010001011: dataB <= 32'b00000111010101011001101011000010;
11'b01010001100: dataB <= 32'b00101100110101000101100001001010;
11'b01010001101: dataB <= 32'b00001010101000110001011010110010;
11'b01010001110: dataB <= 32'b10110101001010001001101000101011;
11'b01010001111: dataB <= 32'b00000100001010010111011011101010;
11'b01010010000: dataB <= 32'b10001011001001010110100011011011;
11'b01010010001: dataB <= 32'b00001100100110101011000100111101;
11'b01010010010: dataB <= 32'b01010110011100100001110011010011;
11'b01010010011: dataB <= 32'b00001001001101100101001010000111;
11'b01010010100: dataB <= 32'b00101101000101010001110110011011;
11'b01010010101: dataB <= 32'b00000101001100000100100010011001;
11'b01010010110: dataB <= 32'b10010001000001101100100110111000;
11'b01010010111: dataB <= 32'b00000101011110010001110101000010;
11'b01010011000: dataB <= 32'b11100000101000110001110000101011;
11'b01010011001: dataB <= 32'b00001101111001100000111110111110;
11'b01010011010: dataB <= 32'b01100001101001001011110011110100;
11'b01010011011: dataB <= 32'b00000101011011000111000101110000;
11'b01010011100: dataB <= 32'b10001111100101100101110100011011;
11'b01010011101: dataB <= 32'b00001011001001101011010101010111;
11'b01010011110: dataB <= 32'b01001010100010101100001011011011;
11'b01010011111: dataB <= 32'b00001010011000011110110101011011;
11'b01010100000: dataB <= 32'b10010111111011000000111101011010;
11'b01010100001: dataB <= 32'b00001000101000100010110101011101;
11'b01010100010: dataB <= 32'b11100011110001011001110111011001;
11'b01010100011: dataB <= 32'b00000110001100011101011101110010;
11'b01010100100: dataB <= 32'b01100111000011011110011011110111;
11'b01010100101: dataB <= 32'b00001110101001110100111010011000;
11'b01010100110: dataB <= 32'b01000010101100111100000011110111;
11'b01010100111: dataB <= 32'b00000100011101001000011000101100;
11'b01010101000: dataB <= 32'b11001001100001010101000010101001;
11'b01010101001: dataB <= 32'b00001010100100101101011101000100;
11'b01010101010: dataB <= 32'b10100100111111110101001101110000;
11'b01010101011: dataB <= 32'b00000111000110011100110010001010;
11'b01010101100: dataB <= 32'b11101111001011001101001011000101;
11'b01010101101: dataB <= 32'b00000010001001001010111011001110;
11'b01010101110: dataB <= 32'b00000000000010010110101000010110;
11'b01010101111: dataB <= 32'b00000000000000000000000000000000;
11'b01010110000: dataB <= 32'b00111000101110111000101110000111;
11'b01010110001: dataB <= 32'b00000100110000101100110100001100;
11'b01010110010: dataB <= 32'b10110101101000101001100101000110;
11'b01010110011: dataB <= 32'b00000010011010010111110011010101;
11'b01010110100: dataB <= 32'b01100100000101100101111000111000;
11'b01010110101: dataB <= 32'b00000000110100010101010001110000;
11'b01010110110: dataB <= 32'b01101100101110000001011000101010;
11'b01010110111: dataB <= 32'b00001001110101110001011000001011;
11'b01010111000: dataB <= 32'b00111011010101001101000111010100;
11'b01010111001: dataB <= 32'b00001010101000111010100000110110;
11'b01010111010: dataB <= 32'b00100000110100001011110100001101;
11'b01010111011: dataB <= 32'b00000100110011111101000001011011;
11'b01010111100: dataB <= 32'b10100101001001111110001010011100;
11'b01010111101: dataB <= 32'b00001100110010010001011101101100;
11'b01010111110: dataB <= 32'b01001110011110010110101100011011;
11'b01010111111: dataB <= 32'b00000001111000101001010101100000;
11'b01011000000: dataB <= 32'b00010000110000110010100110001101;
11'b01011000001: dataB <= 32'b00001111001100010011001010100001;
11'b01011000010: dataB <= 32'b00011111110100111111001100111011;
11'b01011000011: dataB <= 32'b00000100110101000111100001010111;
11'b01011000100: dataB <= 32'b01110010101101100101110111011110;
11'b01011000101: dataB <= 32'b00000101110100110001010111010001;
11'b01011000110: dataB <= 32'b11100010101010000011110101010010;
11'b01011000111: dataB <= 32'b00000001010110111011000101101010;
11'b01011001000: dataB <= 32'b10111101010000011001110000101100;
11'b01011001001: dataB <= 32'b00000110010011001111010101100101;
11'b01011001010: dataB <= 32'b01101100011110110100000100110100;
11'b01011001011: dataB <= 32'b00001110110110110011101110011000;
11'b01011001100: dataB <= 32'b10011010100100110100001110001110;
11'b01011001101: dataB <= 32'b00000000101111100000111010100001;
11'b01011001110: dataB <= 32'b00100010000100010010100011101010;
11'b01011001111: dataB <= 32'b00000001101011010110101000101001;
11'b01011010000: dataB <= 32'b10110110010110111000100100101111;
11'b01011010001: dataB <= 32'b00000100011000011011100001011001;
11'b01011010010: dataB <= 32'b01010110101010001011000110001110;
11'b01011010011: dataB <= 32'b00001011000110100100110001101001;
11'b01011010100: dataB <= 32'b00011011101000010101011100010011;
11'b01011010101: dataB <= 32'b00001001000001011110011110001110;
11'b01011010110: dataB <= 32'b01110001001100001101001000010001;
11'b01011010111: dataB <= 32'b00000001001010101000011101111101;
11'b01011011000: dataB <= 32'b10101110110110001110001110010110;
11'b01011011001: dataB <= 32'b00000110100111100100100010001011;
11'b01011011010: dataB <= 32'b11010100110000001011000100001110;
11'b01011011011: dataB <= 32'b00000011101111100110111100110001;
11'b01011011100: dataB <= 32'b00010100111010111001110010001101;
11'b01011011101: dataB <= 32'b00000100011001101101101110110010;
11'b01011011110: dataB <= 32'b00011001110100011110000101111000;
11'b01011011111: dataB <= 32'b00000010101111110010110110010101;
11'b01011100000: dataB <= 32'b11011100110010101011101110101111;
11'b01011100001: dataB <= 32'b00001010110001110101001101011001;
11'b01011100010: dataB <= 32'b01011010100110110101110101011101;
11'b01011100011: dataB <= 32'b00000100001010101100011101000010;
11'b01011100100: dataB <= 32'b10100100010100110011100101101110;
11'b01011100101: dataB <= 32'b00000101010111101101010001010000;
11'b01011100110: dataB <= 32'b00100101101011010101011101111001;
11'b01011100111: dataB <= 32'b00000011000110100010101010110110;
11'b01011101000: dataB <= 32'b11001111010000111110111001111001;
11'b01011101001: dataB <= 32'b00000110101101100100110111101011;
11'b01011101010: dataB <= 32'b00100010100100111101011101110011;
11'b01011101011: dataB <= 32'b00000110010101010001110100100011;
11'b01011101100: dataB <= 32'b11100001011110010100101100010010;
11'b01011101101: dataB <= 32'b00001111010101111011011101010101;
11'b01011101110: dataB <= 32'b00010100111100111110010101111110;
11'b01011101111: dataB <= 32'b00001100100100011110111111011010;
11'b01011110000: dataB <= 32'b01110100111101111101101010011000;
11'b01011110001: dataB <= 32'b00001101110101100011110000001100;
11'b01011110010: dataB <= 32'b01110011100010111100111101110111;
11'b01011110011: dataB <= 32'b00000100101001101010101011110101;
11'b01011110100: dataB <= 32'b00010001101010000010101101101001;
11'b01011110101: dataB <= 32'b00001100001011011011000001101101;
11'b01011110110: dataB <= 32'b00111101010000011001111101000101;
11'b01011110111: dataB <= 32'b00000100001110011010111010110101;
11'b01011111000: dataB <= 32'b01111000111000111101001100110001;
11'b01011111001: dataB <= 32'b00000110010011101111000101011100;
11'b01011111010: dataB <= 32'b00100000110011001001001011101000;
11'b01011111011: dataB <= 32'b00000100100010011100010100001011;
11'b01011111100: dataB <= 32'b10010111111010000110001011111000;
11'b01011111101: dataB <= 32'b00001110110111001101101110001110;
11'b01011111110: dataB <= 32'b11110001101110100101010100111010;
11'b01011111111: dataB <= 32'b00000010001010101110100110011101;
11'b01100000000: dataB <= 32'b10011110110110100000011000000100;
11'b01100000001: dataB <= 32'b00000011010001011001000101010011;
11'b01100000010: dataB <= 32'b10100100100010100001100010101001;
11'b01100000011: dataB <= 32'b00000100111011011101101011011001;
11'b01100000100: dataB <= 32'b00000000000011010011011011001111;
11'b01100000101: dataB <= 32'b00000000000000000000000000000000;
11'b01100000110: dataB <= 32'b10110010011110001000011011100011;
11'b01100000111: dataB <= 32'b00000101010010101010101100010101;
11'b01100001000: dataB <= 32'b01111011011000010010110011101001;
11'b01100001001: dataB <= 32'b00000100111101100001110111011100;
11'b01100001010: dataB <= 32'b11011000000101111110001010110111;
11'b01100001011: dataB <= 32'b00000010011001011001010101000000;
11'b01100001100: dataB <= 32'b11101000100101100001100111101010;
11'b01100001101: dataB <= 32'b00001010010011110101001000001100;
11'b01100001110: dataB <= 32'b11111100111101011101101000010100;
11'b01100001111: dataB <= 32'b00001001000111110010010001010110;
11'b01100010000: dataB <= 32'b10011110110100001101000011110000;
11'b01100010001: dataB <= 32'b00000101110101111100101101010011;
11'b01100010010: dataB <= 32'b11100111000110010101111100011001;
11'b01100010011: dataB <= 32'b00001100101110010111100101110100;
11'b01100010100: dataB <= 32'b00001000101110110110011110010111;
11'b01100010101: dataB <= 32'b00000011111100101011001100110001;
11'b01100010110: dataB <= 32'b11001110111100101011100101101111;
11'b01100010111: dataB <= 32'b00001101100110010101010010000000;
11'b01100011000: dataB <= 32'b01101001110001101111101110110110;
11'b01100011001: dataB <= 32'b00000110010111010001110001111111;
11'b01100011010: dataB <= 32'b10101100011101111110001001111110;
11'b01100011011: dataB <= 32'b00000111010110110011000110110000;
11'b01100011100: dataB <= 32'b00011110101010000011110101110100;
11'b01100011101: dataB <= 32'b00000011011011111010110001011011;
11'b01100011110: dataB <= 32'b11111100111000001011010000110010;
11'b01100011111: dataB <= 32'b00000111010100010101100001111101;
11'b01100100000: dataB <= 32'b01100100010110110011100101110110;
11'b01100100001: dataB <= 32'b00001111010000111011011001101000;
11'b01100100010: dataB <= 32'b10010110101000111101001101101001;
11'b01100100011: dataB <= 32'b00000001010101100000111010000001;
11'b01100100100: dataB <= 32'b01011000000100001100000011001110;
11'b01100100101: dataB <= 32'b00000001010000010100110000010010;
11'b01100100110: dataB <= 32'b01101100001010001000010100110001;
11'b01100100111: dataB <= 32'b00000110011010100011100000111010;
11'b01100101000: dataB <= 32'b10010100110001111011000110010000;
11'b01100101001: dataB <= 32'b00001001000100100000101101001001;
11'b01100101010: dataB <= 32'b11100011101100101110101100101111;
11'b01100101011: dataB <= 32'b00000110000001011000100010101101;
11'b01100101100: dataB <= 32'b01110010111100100110011000110001;
11'b01100101101: dataB <= 32'b00000000110000100010011010001101;
11'b01100101110: dataB <= 32'b10101100101010101101111111010001;
11'b01100101111: dataB <= 32'b00000101001001011110011110001011;
11'b01100110000: dataB <= 32'b00010010111000001100100100010001;
11'b01100110001: dataB <= 32'b00000100010010100110110100011011;
11'b01100110010: dataB <= 32'b10010101000010011001010010010001;
11'b01100110011: dataB <= 32'b00000110011011110101100010011001;
11'b01100110100: dataB <= 32'b11100101111000111111000111011001;
11'b01100110101: dataB <= 32'b00000011010011101110100110100100;
11'b01100110110: dataB <= 32'b10011000110110100011001101101010;
11'b01100110111: dataB <= 32'b00001010101111110110111101000010;
11'b01100111000: dataB <= 32'b00010110101011001101000111111110;
11'b01100111001: dataB <= 32'b00000011101101100100010100110011;
11'b01100111010: dataB <= 32'b01011100010000110100100101110000;
11'b01100111011: dataB <= 32'b00000110111000101111001000101001;
11'b01100111100: dataB <= 32'b01101101100111011100001111010011;
11'b01100111101: dataB <= 32'b00000001101011011110101011001101;
11'b01100111110: dataB <= 32'b10010101011101100111101011110111;
11'b01100111111: dataB <= 32'b00000110001110100010110011011010;
11'b01101000000: dataB <= 32'b01011110100101010110001110001110;
11'b01101000001: dataB <= 32'b00000111010110011101111000011100;
11'b01101000010: dataB <= 32'b00100111011010011100011100001110;
11'b01101000011: dataB <= 32'b00001111001111111101000101101110;
11'b01101000100: dataB <= 32'b00010111000101100111001000111110;
11'b01101000101: dataB <= 32'b00001010000001011110111111000001;
11'b01101000110: dataB <= 32'b11110000101110001101101011110101;
11'b01101000111: dataB <= 32'b00001110010001101101101100011101;
11'b01101001000: dataB <= 32'b11111001001111000100001110110010;
11'b01101001001: dataB <= 32'b00000011101100100100100111110011;
11'b01101001010: dataB <= 32'b00011011110001110010111100000101;
11'b01101001011: dataB <= 32'b00001010101000011011000101111101;
11'b01101001100: dataB <= 32'b10111100111000001011011011000010;
11'b01101001101: dataB <= 32'b00000100010001011010111110111100;
11'b01101001110: dataB <= 32'b11110110100101010101111100101101;
11'b01101001111: dataB <= 32'b00000111010100101110111001100100;
11'b01101010000: dataB <= 32'b10011110110010100000011010000110;
11'b01101010001: dataB <= 32'b00000010000110010100011000001100;
11'b01101010010: dataB <= 32'b01100011111010011101111101010100;
11'b01101010011: dataB <= 32'b00001111010001011001111010101110;
11'b01101010100: dataB <= 32'b01111001011110101100110111011011;
11'b01101010101: dataB <= 32'b00000001101110101000011010110101;
11'b01101010110: dataB <= 32'b00011100110101110000010110000101;
11'b01101010111: dataB <= 32'b00000011110101011011001101010100;
11'b01101011000: dataB <= 32'b10011110011101111001010010001110;
11'b01101011001: dataB <= 32'b00000111011101100101101010111000;
11'b01101011010: dataB <= 32'b00000000000011001010011010101101;
11'b01101011011: dataB <= 32'b00000000000000000000000000000000;
11'b01101011100: dataB <= 32'b11101010010001100000011001000001;
11'b01101011101: dataB <= 32'b00000101110100100110100100110110;
11'b01101011110: dataB <= 32'b00111101000000001100010010101101;
11'b01101011111: dataB <= 32'b00000111111110101011101111011011;
11'b01101100000: dataB <= 32'b10001110001110011110001011110101;
11'b01101100001: dataB <= 32'b00000100111101011111011000100001;
11'b01101100010: dataB <= 32'b00100010100001001001110110101010;
11'b01101100011: dataB <= 32'b00001011010001110100111000011110;
11'b01101100100: dataB <= 32'b00111010101001110101111001010011;
11'b01101100101: dataB <= 32'b00000111000110100110000101110111;
11'b01101100110: dataB <= 32'b01011100111000100110010100010011;
11'b01101100111: dataB <= 32'b00000110110110110110011001010100;
11'b01101101000: dataB <= 32'b11100111000010101101101101110101;
11'b01101101001: dataB <= 32'b00001100001010011111101001111100;
11'b01101101010: dataB <= 32'b00000111000011001101101111010010;
11'b01101101011: dataB <= 32'b00000110011110101101000000011010;
11'b01101101100: dataB <= 32'b00001111001100101100100101110000;
11'b01101101101: dataB <= 32'b00001011100011011001011001011001;
11'b01101101110: dataB <= 32'b00110011100110010111101111010001;
11'b01101101111: dataB <= 32'b00000111111000011011111010100111;
11'b01101110000: dataB <= 32'b01100110011010011110001100111011;
11'b01101110001: dataB <= 32'b00001000010110110010111010000000;
11'b01101110010: dataB <= 32'b10011010101010000011110110110101;
11'b01101110011: dataB <= 32'b00000101111110110100011101010011;
11'b01101110100: dataB <= 32'b11111010100100001100100001110111;
11'b01101110101: dataB <= 32'b00001000010100011101100110010101;
11'b01101110110: dataB <= 32'b11011100010110100011000111010111;
11'b01101110111: dataB <= 32'b00001111001010111101000101000000;
11'b01101111000: dataB <= 32'b10010010110001010101101100000101;
11'b01101111001: dataB <= 32'b00000010111010011110111001100001;
11'b01101111010: dataB <= 32'b11001100010000010101010011010001;
11'b01101111011: dataB <= 32'b00000010010101010010111100001011;
11'b01101111100: dataB <= 32'b00100000000101100000010101110011;
11'b01101111101: dataB <= 32'b00001000011011101001011100110011;
11'b01101111110: dataB <= 32'b01010010111101110011000110010001;
11'b01101111111: dataB <= 32'b00000110100100011110101100110010;
11'b01110000000: dataB <= 32'b01101011100101010111011100001100;
11'b01110000001: dataB <= 32'b00000011100011010010101010111101;
11'b01110000010: dataB <= 32'b00110000110001001111011000110001;
11'b01110000011: dataB <= 32'b00000001010101011010011110011101;
11'b01110000100: dataB <= 32'b01100110100010111101011110101011;
11'b01110000101: dataB <= 32'b00000011101011011000100010000011;
11'b01110000110: dataB <= 32'b01010011000100011101110100110100;
11'b01110000111: dataB <= 32'b00000100110101100100110000011100;
11'b01110001000: dataB <= 32'b10010101001001111001000010110110;
11'b01110001001: dataB <= 32'b00001000111011111011001101111001;
11'b01110001010: dataB <= 32'b01101111110001100111101001011000;
11'b01110001011: dataB <= 32'b00000011110110101000011110101100;
11'b01110001100: dataB <= 32'b01011000111010011010111100000110;
11'b01110001101: dataB <= 32'b00001010101101110100101100110011;
11'b01110001110: dataB <= 32'b00010010110011010100001010111101;
11'b01110001111: dataB <= 32'b00000011010001011100010100110100;
11'b01110010000: dataB <= 32'b10010100011001000101010110010010;
11'b01110010001: dataB <= 32'b00001000111001101110111100010010;
11'b01110010010: dataB <= 32'b01110011011011010011001111001110;
11'b01110010011: dataB <= 32'b00000001010000011010101011011100;
11'b01110010100: dataB <= 32'b10011011100110010111101100110011;
11'b01110010101: dataB <= 32'b00000110001111100000110011000001;
11'b01110010110: dataB <= 32'b01011000101001110110011101101010;
11'b01110010111: dataB <= 32'b00001000110110101001111000100101;
11'b01110011000: dataB <= 32'b01101011010010011100001011101011;
11'b01110011001: dataB <= 32'b00001110101001111100110010001110;
11'b01110011010: dataB <= 32'b10011001001110001111001011011101;
11'b01110011011: dataB <= 32'b00000111100001011110111110011000;
11'b01110011100: dataB <= 32'b11101100100010011101001100110010;
11'b01110011101: dataB <= 32'b00001110001100110101100000110110;
11'b01110011110: dataB <= 32'b01111000111011000011001110101101;
11'b01110011111: dataB <= 32'b00000011001111100000100011101010;
11'b01110100000: dataB <= 32'b00100101110001100011001001100010;
11'b01110100001: dataB <= 32'b00001001000110011101001010001101;
11'b01110100010: dataB <= 32'b11111010100000001100101000000001;
11'b01110100011: dataB <= 32'b00000100110100011011000010111011;
11'b01110100100: dataB <= 32'b00110000010101101110011011101010;
11'b01110100101: dataB <= 32'b00001000010100101100101101110101;
11'b01110100110: dataB <= 32'b11011100110101110000011000000101;
11'b01110100111: dataB <= 32'b00000000101011001110100100011101;
11'b01110101000: dataB <= 32'b10101101110110110101011101110000;
11'b01110101001: dataB <= 32'b00001111001011100011111011000101;
11'b01110101010: dataB <= 32'b10111101001010110100001001111011;
11'b01110101011: dataB <= 32'b00000001110011100000010110111100;
11'b01110101100: dataB <= 32'b10011010111001000000100100000111;
11'b01110101101: dataB <= 32'b00000101011000011101001101010100;
11'b01110101110: dataB <= 32'b01011000100001011001100010010011;
11'b01110101111: dataB <= 32'b00001001111101101101100010001000;
11'b01110110000: dataB <= 32'b00000000000010110001101010001011;
11'b01110110001: dataB <= 32'b00000000000000000000000000000000;
11'b01110110010: dataB <= 32'b10100000001000110001000110000001;
11'b01110110011: dataB <= 32'b00000110110101100000100001011111;
11'b01110110100: dataB <= 32'b00111100101000011101100010110001;
11'b01110110101: dataB <= 32'b00001010111110110011100111001010;
11'b01110110110: dataB <= 32'b00000110011110101101101100010001;
11'b01110110111: dataB <= 32'b00000111111110100011011000001011;
11'b01110111000: dataB <= 32'b00011100100000110010110101101100;
11'b01110111001: dataB <= 32'b00001011001111110010101000111111;
11'b01110111010: dataB <= 32'b11110100010110001101111001110010;
11'b01110111011: dataB <= 32'b00000101100111011100000110011110;
11'b01110111100: dataB <= 32'b11011100111001001111010101010110;
11'b01110111101: dataB <= 32'b00001000010111101100001001011100;
11'b01110111110: dataB <= 32'b11100110111010111100111110110000;
11'b01110111111: dataB <= 32'b00001010100111101001100110001100;
11'b01111000000: dataB <= 32'b10001001010011010100101110101100;
11'b01111000001: dataB <= 32'b00001001011110101100111000001011;
11'b01111000010: dataB <= 32'b11010011010100111101100110010010;
11'b01111000011: dataB <= 32'b00001000100001011111011100111001;
11'b01111000100: dataB <= 32'b01111001010111000111001111001011;
11'b01111000101: dataB <= 32'b00001001010111100111111011001110;
11'b01111000110: dataB <= 32'b01011110010110101101101110110111;
11'b01111000111: dataB <= 32'b00001001010101110000101001010000;
11'b01111001000: dataB <= 32'b00010110110010000011110111110110;
11'b01111001001: dataB <= 32'b00001000011110101100010001010100;
11'b01111001010: dataB <= 32'b10110010010000011110000011111100;
11'b01111001011: dataB <= 32'b00001001010100100101100110100101;
11'b01111001100: dataB <= 32'b11010100011010011010101000110111;
11'b01111001101: dataB <= 32'b00001101100101111100101100011001;
11'b01111001110: dataB <= 32'b00010000111101101110001001100011;
11'b01111001111: dataB <= 32'b00000101011101011110111001001010;
11'b01111010000: dataB <= 32'b01000100100000101110100011110101;
11'b01111010001: dataB <= 32'b00000011011001010011000100001101;
11'b01111010010: dataB <= 32'b00010100000100110001000110010101;
11'b01111010011: dataB <= 32'b00001010111010101111010100101100;
11'b01111010100: dataB <= 32'b01010011000101101011010110110010;
11'b01111010101: dataB <= 32'b00000100100110011010110000101011;
11'b01111010110: dataB <= 32'b01110001011010000111101011001001;
11'b01111010111: dataB <= 32'b00000001100111010000110111000100;
11'b01111011000: dataB <= 32'b10101100100101111111101000110000;
11'b01111011001: dataB <= 32'b00000010111010010100100010100100;
11'b01111011010: dataB <= 32'b01100000011111000100011101000110;
11'b01111011011: dataB <= 32'b00000011001111010010101001111011;
11'b01111011100: dataB <= 32'b01010101001100111111000101110110;
11'b01111011101: dataB <= 32'b00000110010111100000110000100101;
11'b01111011110: dataB <= 32'b10011001010001010001010100011001;
11'b01111011111: dataB <= 32'b00001011011010111010111001011001;
11'b01111100000: dataB <= 32'b11110111100010010111101010110111;
11'b01111100001: dataB <= 32'b00000101111001100000010110101011;
11'b01111100010: dataB <= 32'b01010111000010001010101010000011;
11'b01111100011: dataB <= 32'b00001001101011101110011100110100;
11'b01111100100: dataB <= 32'b00010000111111001011001101011010;
11'b01111100101: dataB <= 32'b00000011110100010100011000110101;
11'b01111100110: dataB <= 32'b00001110100101011110000110110011;
11'b01111100111: dataB <= 32'b00001010011000101100110000001100;
11'b01111101000: dataB <= 32'b01110101001011000010001110101000;
11'b01111101001: dataB <= 32'b00000001110101010110110011010011;
11'b01111101010: dataB <= 32'b11100011100110111111001101001111;
11'b01111101011: dataB <= 32'b00000110010001011100110010100000;
11'b01111101100: dataB <= 32'b01010100101110010110011100000110;
11'b01111101101: dataB <= 32'b00001001110101110011101100111110;
11'b01111101110: dataB <= 32'b00101101001010011011101010101000;
11'b01111101111: dataB <= 32'b00001101000101110110011010100110;
11'b01111110000: dataB <= 32'b10011101010010101110111101111001;
11'b01111110001: dataB <= 32'b00000100100010011110111101101000;
11'b01111110010: dataB <= 32'b10100100011010101100111100101110;
11'b01111110011: dataB <= 32'b00001100100111111001001101100111;
11'b01111110100: dataB <= 32'b01110110101010110010101101101000;
11'b01111110101: dataB <= 32'b00000011110011011010100111010001;
11'b01111110110: dataB <= 32'b11101111101001011011100111000010;
11'b01111110111: dataB <= 32'b00000111000110011111001010011100;
11'b01111111000: dataB <= 32'b00110010010000011110000101000001;
11'b01111111001: dataB <= 32'b00000101110110011011000110110011;
11'b01111111010: dataB <= 32'b01100110001110001110011010000111;
11'b01111111011: dataB <= 32'b00001001010100101000100110000101;
11'b01111111100: dataB <= 32'b00011010111001000000100101100110;
11'b01111111101: dataB <= 32'b00000000110000001010110000111111;
11'b01111111110: dataB <= 32'b11110111100110111100101101001100;
11'b01111111111: dataB <= 32'b00001101100110101111110111010100;
11'b10000000000: dataB <= 32'b11111010110010110011101011111001;
11'b10000000001: dataB <= 32'b00000011011000011000011011000011;
11'b10000000010: dataB <= 32'b00011010111100100001100010101010;
11'b10000000011: dataB <= 32'b00000111011001100001010001100101;
11'b10000000100: dataB <= 32'b01010010101001000010000011010111;
11'b10000000101: dataB <= 32'b00001100011010110011010101011000;
11'b10000000110: dataB <= 32'b00000000000010010001011001001010;
11'b10000000111: dataB <= 32'b00000000000000000000000000000000;
11'b10000001000: dataB <= 32'b00000100111100100110010000110011;
11'b10000001001: dataB <= 32'b00001010110010010000111111110101;
11'b10000001010: dataB <= 32'b10010100000110110111001000111010;
11'b10000001011: dataB <= 32'b00001111001010110010011001000001;
11'b10000001100: dataB <= 32'b10001111110010110010101000100111;
11'b10000001101: dataB <= 32'b00001111010000101100111001100111;
11'b10000001110: dataB <= 32'b00010001000101011110010110010100;
11'b10000001111: dataB <= 32'b00000111101001010100011011100110;
11'b10000010000: dataB <= 32'b00001010010110111011101001001100;
11'b10000010001: dataB <= 32'b00000011110100000011000111011011;
11'b10000010010: dataB <= 32'b00011101000111101101101011010101;
11'b10000010011: dataB <= 32'b00001011101111000100100110011101;
11'b10000010100: dataB <= 32'b10011100110010011010001000000010;
11'b10000010101: dataB <= 32'b00000011101010110010101110011011;
11'b10000010110: dataB <= 32'b10101001101110010001010110000010;
11'b10000010111: dataB <= 32'b00001111001101011100100101110111;
11'b10000011000: dataB <= 32'b00101011011010110110001001010011;
11'b10000011001: dataB <= 32'b00000000101110101111000000111110;
11'b10000011010: dataB <= 32'b10101010001111100001110101100001;
11'b10000011011: dataB <= 32'b00001011101101111100110011001001;
11'b10000011100: dataB <= 32'b01001011000010110010101011100010;
11'b10000011101: dataB <= 32'b00001010101101010100011100001101;
11'b10000011110: dataB <= 32'b01011001010001111011111011010000;
11'b10000011111: dataB <= 32'b00001111001111001000100110000101;
11'b10000100000: dataB <= 32'b11001000011011000111001110011000;
11'b10000100001: dataB <= 32'b00001010001101110010110110110010;
11'b10000100010: dataB <= 32'b00001101010101010011001011101110;
11'b10000100011: dataB <= 32'b00000010100100010110000100111111;
11'b10000100100: dataB <= 32'b10011111011111000100100001101100;
11'b10000100101: dataB <= 32'b00001110110101011101000001000101;
11'b10000100110: dataB <= 32'b10010001110111010110101010111000;
11'b10000100111: dataB <= 32'b00001100111001100011011010101111;
11'b10000101000: dataB <= 32'b10000011010100100110011010110011;
11'b10000101001: dataB <= 32'b00001101001010101010100010000110;
11'b10000101010: dataB <= 32'b10100011011001101100101001010010;
11'b10000101011: dataB <= 32'b00000011010110011001001001101110;
11'b10000101100: dataB <= 32'b11101100011111110011110100101001;
11'b10000101101: dataB <= 32'b00000011111100011011011110001001;
11'b10000101110: dataB <= 32'b11010010100111110100001000001110;
11'b10000101111: dataB <= 32'b00001101011010010001010110010010;
11'b10000110000: dataB <= 32'b00001110111110001001110011000101;
11'b10000110001: dataB <= 32'b00000111111001010101011001101100;
11'b10000110010: dataB <= 32'b11100111010111100110001011010100;
11'b10000110011: dataB <= 32'b00001011110011011000111110101110;
11'b10000110100: dataB <= 32'b00101001001100101101011100110111;
11'b10000110101: dataB <= 32'b00001101001001011100001000110101;
11'b10000110110: dataB <= 32'b10110000010011110011011011101010;
11'b10000110111: dataB <= 32'b00001100110100001010111101111010;
11'b10000111000: dataB <= 32'b01100001010001010011100001101011;
11'b10000111001: dataB <= 32'b00000101101100001110100010001110;
11'b10000111010: dataB <= 32'b01011111011101100001101101000101;
11'b10000111011: dataB <= 32'b00001010011000001101010110100110;
11'b10000111100: dataB <= 32'b10010011100011000101001001110010;
11'b10000111101: dataB <= 32'b00001100001011011000100110000111;
11'b10000111110: dataB <= 32'b01100100010101000001110100000010;
11'b10000111111: dataB <= 32'b00001010111100011001010001101001;
11'b10001000000: dataB <= 32'b11110010111011100010000111100101;
11'b10001000001: dataB <= 32'b00001000110011011001000100011010;
11'b10001000010: dataB <= 32'b00010111010111001011010011000111;
11'b10001000011: dataB <= 32'b00001010101100110110011011001110;
11'b10001000100: dataB <= 32'b11100100100101110011000100001010;
11'b10001000101: dataB <= 32'b00000010100101001100010011000010;
11'b10001000110: dataB <= 32'b10101001000111011010101100100100;
11'b10001000111: dataB <= 32'b00000001010110011111000000010100;
11'b10001001000: dataB <= 32'b11001100110110011010100111000110;
11'b10001001001: dataB <= 32'b00000011100110100110001111110100;
11'b10001001010: dataB <= 32'b01010100010001010010010100000100;
11'b10001001011: dataB <= 32'b00001001111000010011001000101001;
11'b10001001100: dataB <= 32'b00110100100001110101000001010001;
11'b10001001101: dataB <= 32'b00000011010001100101000010011011;
11'b10001001110: dataB <= 32'b01001000011011000111000000110101;
11'b10001001111: dataB <= 32'b00001011010100100011001001100010;
11'b10001010000: dataB <= 32'b11000110110011001011100011101011;
11'b10001010001: dataB <= 32'b00001010001101010010101110101011;
11'b10001010010: dataB <= 32'b00011101001000010101110011010100;
11'b10001010011: dataB <= 32'b00001000011110011001101011100110;
11'b10001010100: dataB <= 32'b01110010010010010010000110000101;
11'b10001010101: dataB <= 32'b00000011000100111010100010011001;
11'b10001010110: dataB <= 32'b11011000001001110010011100101000;
11'b10001010111: dataB <= 32'b00001100011001001101001101111001;
11'b10001011000: dataB <= 32'b11011111001000110110110101011010;
11'b10001011001: dataB <= 32'b00001100110001101000111110100100;
11'b10001011010: dataB <= 32'b00010101011001000101111011111001;
11'b10001011011: dataB <= 32'b00001101000111101010011000001101;
11'b10001011100: dataB <= 32'b00000000000000101011010101001101;
11'b10001011101: dataB <= 32'b00000000000000000000000000000000;
11'b10001011110: dataB <= 32'b01001000101000001100110000101101;
11'b10001011111: dataB <= 32'b00001010010100010010110011011110;
11'b10001100000: dataB <= 32'b00100000000110001111100110111010;
11'b10001100001: dataB <= 32'b00001111010000110110101001100001;
11'b10001100010: dataB <= 32'b11000111100011000011001010101000;
11'b10001100011: dataB <= 32'b00001110110110101101000000110110;
11'b10001100100: dataB <= 32'b00010000111000111101100101010010;
11'b10001100101: dataB <= 32'b00001000101001011100010111000111;
11'b10001100110: dataB <= 32'b01010100001010111100011001101101;
11'b10001100111: dataB <= 32'b00000011010001000010110011100100;
11'b10001101000: dataB <= 32'b01011101000111001110111001110111;
11'b10001101001: dataB <= 32'b00001011010010001100010010001101;
11'b10001101010: dataB <= 32'b00100000110010110010101010100100;
11'b10001101011: dataB <= 32'b00000101000111110101000010011100;
11'b10001101100: dataB <= 32'b00100001110010110001101001000001;
11'b10001101101: dataB <= 32'b00001111010011100000100101000111;
11'b10001101110: dataB <= 32'b00100111100010010110101000010100;
11'b10001101111: dataB <= 32'b00000001101000101101001100100101;
11'b10001110000: dataB <= 32'b11110010011011110011011000100001;
11'b10001110001: dataB <= 32'b00001100010000111101001011100010;
11'b10001110010: dataB <= 32'b11001100110011000011001101100110;
11'b10001110011: dataB <= 32'b00001011001111011100011000001011;
11'b10001110100: dataB <= 32'b01010101001001111011111010110010;
11'b10001110101: dataB <= 32'b00001111010100001110010101110101;
11'b10001110110: dataB <= 32'b01010010001010010111101011111100;
11'b10001110111: dataB <= 32'b00001010001111110011000110111011;
11'b10001111000: dataB <= 32'b11001011000101100010111011110001;
11'b10001111001: dataB <= 32'b00000101000001100010000100011101;
11'b10001111010: dataB <= 32'b11011001011010110101010010100111;
11'b10001111011: dataB <= 32'b00001101011010011101000000110100;
11'b10001111100: dataB <= 32'b10001001100110101111011000111001;
11'b10001111101: dataB <= 32'b00001010111011011111011001111111;
11'b10001111110: dataB <= 32'b01000010111100001100111001110100;
11'b10001111111: dataB <= 32'b00001101101111101110101101100110;
11'b10010000000: dataB <= 32'b01011111011001100100011000110011;
11'b10010000001: dataB <= 32'b00000010010010010111000001001110;
11'b10010000010: dataB <= 32'b00110010101011101101010110000111;
11'b10010000011: dataB <= 32'b00000001111000010101011010101010;
11'b10010000100: dataB <= 32'b00011000011111101101101000101110;
11'b10010000101: dataB <= 32'b00001010111101001111001010100011;
11'b10010000110: dataB <= 32'b11010000110010101010000101100010;
11'b10010000111: dataB <= 32'b00000101111000010001001101101011;
11'b10010001000: dataB <= 32'b00100011011010111111001010010110;
11'b10010001001: dataB <= 32'b00001010110110011000110110001111;
11'b10010001010: dataB <= 32'b00100101010100100100001011011010;
11'b10010001011: dataB <= 32'b00001101101110100110001000110100;
11'b10010001100: dataB <= 32'b10111000100011110100111100001101;
11'b10010001101: dataB <= 32'b00001011011000001110101110001010;
11'b10010001110: dataB <= 32'b01011101001101011011000011000111;
11'b10010001111: dataB <= 32'b00000110101010010110010101101110;
11'b10010010000: dataB <= 32'b01011001011010000001011110101010;
11'b10010010001: dataB <= 32'b00001000111001001011000110000110;
11'b10010010010: dataB <= 32'b01001101010110101101111001010011;
11'b10010010011: dataB <= 32'b00001100101110011110100001010111;
11'b10010010100: dataB <= 32'b00101100011001100001010111000001;
11'b10010010101: dataB <= 32'b00001000011101010101001010001001;
11'b10010010110: dataB <= 32'b11110011001011110011011001100110;
11'b10010010111: dataB <= 32'b00000111110011011000111100110001;
11'b10010011000: dataB <= 32'b11010101001111001100010101000100;
11'b10010011001: dataB <= 32'b00001011001110111100101110101110;
11'b10010011010: dataB <= 32'b10101000101010000011000101101000;
11'b10010011011: dataB <= 32'b00000100100010011000000111001011;
11'b10010011100: dataB <= 32'b00100111001111100011101110101001;
11'b10010011101: dataB <= 32'b00000000110000011111000000010011;
11'b10010011110: dataB <= 32'b01010000100110100011001001000110;
11'b10010011111: dataB <= 32'b00000110000011110000010111011110;
11'b10010100000: dataB <= 32'b10011100001101100001110110100010;
11'b10010100001: dataB <= 32'b00000111111001010000111101001000;
11'b10010100010: dataB <= 32'b10111000110101100100110001001100;
11'b10010100011: dataB <= 32'b00000011001101100101000110100011;
11'b10010100100: dataB <= 32'b00010000001010010111100000101111;
11'b10010100101: dataB <= 32'b00001010010110100001001001111010;
11'b10010100110: dataB <= 32'b01001010011111001100100101001000;
11'b10010100111: dataB <= 32'b00001010001111010110100110100100;
11'b10010101000: dataB <= 32'b00011011000100001100010010101111;
11'b10010101001: dataB <= 32'b00000101111110010011100010111111;
11'b10010101010: dataB <= 32'b11111010100110101010011000000100;
11'b10010101011: dataB <= 32'b00000101100001111100111010110001;
11'b10010101100: dataB <= 32'b00100100000110000010011101101100;
11'b10010101101: dataB <= 32'b00001001111100001010111110010010;
11'b10010101110: dataB <= 32'b01011101001000010101110011110111;
11'b10010101111: dataB <= 32'b00001100010101100111000110010101;
11'b10010110000: dataB <= 32'b10010001001100110101001001111011;
11'b10010110001: dataB <= 32'b00001110101100110000100100001011;
11'b10010110010: dataB <= 32'b00000000000000110010010101101011;
11'b10010110011: dataB <= 32'b00000000000000000000000000000000;
11'b10010110100: dataB <= 32'b01001110011000001011100001101000;
11'b10010110101: dataB <= 32'b00001001010101010110101010110111;
11'b10010110110: dataB <= 32'b00101100001001011111010100111000;
11'b10010110111: dataB <= 32'b00001110110110111010111110001001;
11'b10010111000: dataB <= 32'b11000011001111000100001011101010;
11'b10010111001: dataB <= 32'b00001100111011101011001100011101;
11'b10010111010: dataB <= 32'b10010010101100110100110101010000;
11'b10010111011: dataB <= 32'b00001001101011100100010110011111;
11'b10010111100: dataB <= 32'b01011110000110110101001010001111;
11'b10010111101: dataB <= 32'b00000011101101001000011011011101;
11'b10010111110: dataB <= 32'b01011011000010100111101000011000;
11'b10010111111: dataB <= 32'b00001010110100010110000101110101;
11'b10011000000: dataB <= 32'b01100010110010111011011100100111;
11'b10011000001: dataB <= 32'b00000111000110110011010010011100;
11'b10011000010: dataB <= 32'b01010111101111001010011011100011;
11'b10011000011: dataB <= 32'b00001110011000100110101000100110;
11'b10011000100: dataB <= 32'b11011111100001110110100111110100;
11'b10011000101: dataB <= 32'b00000011000100101001010100011011;
11'b10011000110: dataB <= 32'b00111000101111110100101011000010;
11'b10011000111: dataB <= 32'b00001011110011111001011111101100;
11'b10011001000: dataB <= 32'b01001110100111000100001111001100;
11'b10011001001: dataB <= 32'b00001011010001100010011000010010;
11'b10011001010: dataB <= 32'b00010101000001111011111010010100;
11'b10011001011: dataB <= 32'b00001101111001011000001001100101;
11'b10011001100: dataB <= 32'b00011100000101101111101001011110;
11'b10011001101: dataB <= 32'b00001010010001110001010110111100;
11'b10011001110: dataB <= 32'b10001010110101110010011011010100;
11'b10011001111: dataB <= 32'b00001000000001101100001000001100;
11'b10011010000: dataB <= 32'b11010101010010100110000100100100;
11'b10011010001: dataB <= 32'b00001010111101011100111100110011;
11'b10011010010: dataB <= 32'b01000011001110000111100111011001;
11'b10011010011: dataB <= 32'b00001000011101011001010101001111;
11'b10011010100: dataB <= 32'b00000100100100001011101000110110;
11'b10011010101: dataB <= 32'b00001101010011110000111001001110;
11'b10011010110: dataB <= 32'b10011001010101100100001000010011;
11'b10011010111: dataB <= 32'b00000010001101010110111100110101;
11'b10011011000: dataB <= 32'b10110110111011010110100111100110;
11'b10011011001: dataB <= 32'b00000000110011010001001110111010;
11'b10011011010: dataB <= 32'b10011110011011001110111000101110;
11'b10011011011: dataB <= 32'b00001000011110001100111010101011;
11'b10011011100: dataB <= 32'b10010100100110111010101000100001;
11'b10011011101: dataB <= 32'b00000100110101001111000001110011;
11'b10011011110: dataB <= 32'b00011101011010010111101000110111;
11'b10011011111: dataB <= 32'b00001001010111011010110001100111;
11'b10011100000: dataB <= 32'b00100001010100101011001000111011;
11'b10011100001: dataB <= 32'b00001101110011110000010100110011;
11'b10011100010: dataB <= 32'b11111100110111100110001100110001;
11'b10011100011: dataB <= 32'b00001001111001010010100010011010;
11'b10011100100: dataB <= 32'b11011011001101100010110101000100;
11'b10011100101: dataB <= 32'b00000111101010011110010001010101;
11'b10011100110: dataB <= 32'b01010101010010100001101111010000;
11'b10011100111: dataB <= 32'b00000110111000001010110101100110;
11'b10011101000: dataB <= 32'b10001001000110010110011000010100;
11'b10011101001: dataB <= 32'b00001100010010100100100000101110;
11'b10011101010: dataB <= 32'b10110010100110000001001001100001;
11'b10011101011: dataB <= 32'b00000101111100010101000010101001;
11'b10011101100: dataB <= 32'b00101111010111110100111011101000;
11'b10011101101: dataB <= 32'b00000111010011011000111001010001;
11'b10011101110: dataB <= 32'b00010011000011000101010111000011;
11'b10011101111: dataB <= 32'b00001011010001111101000110001111;
11'b10011110000: dataB <= 32'b10101100110010001011000111000111;
11'b10011110001: dataB <= 32'b00000111100001100010000111000100;
11'b10011110010: dataB <= 32'b11100011010011100100111111001110;
11'b10011110011: dataB <= 32'b00000000101011011111000000100001;
11'b10011110100: dataB <= 32'b00010110011110110011101010101000;
11'b10011110101: dataB <= 32'b00001000100011110110100110111111;
11'b10011110110: dataB <= 32'b01100110001110000001111001000010;
11'b10011110111: dataB <= 32'b00000110011000010010110101111000;
11'b10011111000: dataB <= 32'b00111001001001011100010010100111;
11'b10011111001: dataB <= 32'b00000100001010100011001010100100;
11'b10011111010: dataB <= 32'b00011100000101101111100001001001;
11'b10011111011: dataB <= 32'b00001000110111011111001010010010;
11'b10011111100: dataB <= 32'b11010010010010111101010110100110;
11'b10011111101: dataB <= 32'b00001010010001011100100010011100;
11'b10011111110: dataB <= 32'b10011001000000001010110011001011;
11'b10011111111: dataB <= 32'b00000011011011001101010110010111;
11'b10100000000: dataB <= 32'b10111100111010111011001010000101;
11'b10100000001: dataB <= 32'b00001000100001111101001111001010;
11'b10100000010: dataB <= 32'b01101110001110011010101101110001;
11'b10100000011: dataB <= 32'b00000111011100001100101110101010;
11'b10100000100: dataB <= 32'b01011011000100001100010010110011;
11'b10100000101: dataB <= 32'b00001010111000100111001010000101;
11'b10100000110: dataB <= 32'b00001111000000101100000111011011;
11'b10100000111: dataB <= 32'b00001110110001110100110100010010;
11'b10100001000: dataB <= 32'b00000000000001001001100110101010;
11'b10100001001: dataB <= 32'b00000000000000000000000000000000;
11'b10100001010: dataB <= 32'b10010110001100010010000011100011;
11'b10100001011: dataB <= 32'b00001000010110011010100110000111;
11'b10100001100: dataB <= 32'b01110100010100110110100011010101;
11'b10100001101: dataB <= 32'b00001101011011111001010010110001;
11'b10100001110: dataB <= 32'b01000010110110111100111100001110;
11'b10100001111: dataB <= 32'b00001010011110101001010100001100;
11'b10100010000: dataB <= 32'b10010110100100101011110101001110;
11'b10100010001: dataB <= 32'b00001010101100101100011101101111;
11'b10100010010: dataB <= 32'b01101010001010100101101010010001;
11'b10100010011: dataB <= 32'b00000100001010010000001011000110;
11'b10100010100: dataB <= 32'b00011010111101111111100110110111;
11'b10100010101: dataB <= 32'b00001001110110100000000101100101;
11'b10100010110: dataB <= 32'b10100100110111000100001110001011;
11'b10100010111: dataB <= 32'b00001001000110101111011110010100;
11'b10100011000: dataB <= 32'b11001111100011010011011101100111;
11'b10100011001: dataB <= 32'b00001100011100101010101100001100;
11'b10100011010: dataB <= 32'b11011001011101010110010110110011;
11'b10100011011: dataB <= 32'b00000110000001100101011000100010;
11'b10100011100: dataB <= 32'b01111011000011100110001101100110;
11'b10100011101: dataB <= 32'b00001010110110110001110011100101;
11'b10100011110: dataB <= 32'b01010110011010111100111111010001;
11'b10100011111: dataB <= 32'b00001010010100101010011100101001;
11'b10100100000: dataB <= 32'b10010100111001111011111001010101;
11'b10100100001: dataB <= 32'b00001011011101100010001001011100;
11'b10100100010: dataB <= 32'b11101000000100111111000110011110;
11'b10100100011: dataB <= 32'b00001001110011101011100010110100;
11'b10100100100: dataB <= 32'b00001110100110000010011010010110;
11'b10100100101: dataB <= 32'b00001011000010110110011000001011;
11'b10100100110: dataB <= 32'b11010011001010000110010111000011;
11'b10100100111: dataB <= 32'b00000111111110011100111100110010;
11'b10100101000: dataB <= 32'b10000010111001010111010101011000;
11'b10100101001: dataB <= 32'b00000101111100010101010000100110;
11'b10100101010: dataB <= 32'b00001010010000010010000111110110;
11'b10100101011: dataB <= 32'b00001100010111110001001000110101;
11'b10100101100: dataB <= 32'b10010101010001100011100111010011;
11'b10100101101: dataB <= 32'b00000011001001011000110100101100;
11'b10100101110: dataB <= 32'b10110101001010101111011001100111;
11'b10100101111: dataB <= 32'b00000000101101001111000011000011;
11'b10100110000: dataB <= 32'b00100110011110100111101000101111;
11'b10100110001: dataB <= 32'b00000101011101001110101110101100;
11'b10100110010: dataB <= 32'b10011010100011000011101011000011;
11'b10100110011: dataB <= 32'b00000011110010010000110101110011;
11'b10100110100: dataB <= 32'b01011001010101100111100111010111;
11'b10100110101: dataB <= 32'b00000111111000011110110000111110;
11'b10100110110: dataB <= 32'b01011101010100111010000110111011;
11'b10100110111: dataB <= 32'b00001100110111110110100101000010;
11'b10100111000: dataB <= 32'b01111011001111000111001100010100;
11'b10100111001: dataB <= 32'b00000111111010011010011010100011;
11'b10100111010: dataB <= 32'b00011001000101110010100111100010;
11'b10100111011: dataB <= 32'b00001000101010100110010100111101;
11'b10100111100: dataB <= 32'b11010011001010111010011110110101;
11'b10100111101: dataB <= 32'b00000101010111001110100101001101;
11'b10100111110: dataB <= 32'b01001010110101110110010111010100;
11'b10100111111: dataB <= 32'b00001011110101101000100100010101;
11'b10101000000: dataB <= 32'b01110100110110101001011100100100;
11'b10101000001: dataB <= 32'b00000011011001010100111011000010;
11'b10101000010: dataB <= 32'b10101001100011011110001100101100;
11'b10101000011: dataB <= 32'b00000110110010011010110101111000;
11'b10101000100: dataB <= 32'b11010010111010101110001001100100;
11'b10101000101: dataB <= 32'b00001010110011111011011101100110;
11'b10101000110: dataB <= 32'b01101110111110010011011001000111;
11'b10101000111: dataB <= 32'b00001010100001101110001010111101;
11'b10101001000: dataB <= 32'b00011111010111001110001111010100;
11'b10101001001: dataB <= 32'b00000010000110011111000001000001;
11'b10101001010: dataB <= 32'b10011110010110110100001100001011;
11'b10101001011: dataB <= 32'b00001010100100111000111010001111;
11'b10101001100: dataB <= 32'b01110000011010011010001011100100;
11'b10101001101: dataB <= 32'b00000100110110010100101010101000;
11'b10101001110: dataB <= 32'b10110101011101010011110100100100;
11'b10101001111: dataB <= 32'b00000101100111100001001010100100;
11'b10101010000: dataB <= 32'b01101000000100111111000010100101;
11'b10101010001: dataB <= 32'b00000111010111011101001010100010;
11'b10101010010: dataB <= 32'b00011100001110100110001000100110;
11'b10101010011: dataB <= 32'b00001001110011100010100010001101;
11'b10101010100: dataB <= 32'b10011000111100100001100100001000;
11'b10101010101: dataB <= 32'b00000001010110001011000101100111;
11'b10101010110: dataB <= 32'b10111101010011000011111100001000;
11'b10101010111: dataB <= 32'b00001011100010110111100111010011;
11'b10101011000: dataB <= 32'b00110110011110101010111101010110;
11'b10101011001: dataB <= 32'b00000101011011010010100010111011;
11'b10101011010: dataB <= 32'b01011011000000001010110010001111;
11'b10101011011: dataB <= 32'b00001000111001100011001101110101;
11'b10101011100: dataB <= 32'b00010000110100110010110100111010;
11'b10101011101: dataB <= 32'b00001101110110110101000100110001;
11'b10101011110: dataB <= 32'b00000000000001101001010111101001;
11'b10101011111: dataB <= 32'b00000000000000000000000000000000;
endcase
end
assign doA = dataA;
assign doB = dataB;
endmodule
